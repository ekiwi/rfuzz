module Sodor5Stage(
  input          metaReset,
  input          clock,
  input          reset,
  input          io_imem_req_ready,
  output         io_imem_req_valid,
  output [31:0]  io_imem_req_bits_addr,
  output [31:0]  io_imem_req_bits_data,
  output         io_imem_req_bits_fcn,
  output [2:0]   io_imem_req_bits_typ,
  input          io_imem_resp_valid,
  input  [31:0]  io_imem_resp_bits_data,
  input          io_reset,
  output         assert_out,
  output [791:0] auto_cover_out
);
  wire  core_metaReset; // @[top.scala 21:26]
  wire  core_clock; // @[top.scala 21:26]
  wire  core_reset; // @[top.scala 21:26]
  wire [31:0] core_io_imem_req_bits_addr; // @[top.scala 21:26]
  wire  core_io_imem_resp_valid; // @[top.scala 21:26]
  wire [31:0] core_io_imem_resp_bits_data; // @[top.scala 21:26]
  wire  core_io_dmem_req_valid; // @[top.scala 21:26]
  wire [31:0] core_io_dmem_req_bits_addr; // @[top.scala 21:26]
  wire [31:0] core_io_dmem_req_bits_data; // @[top.scala 21:26]
  wire  core_io_dmem_req_bits_fcn; // @[top.scala 21:26]
  wire [2:0] core_io_dmem_req_bits_typ; // @[top.scala 21:26]
  wire  core_io_dmem_resp_valid; // @[top.scala 21:26]
  wire [31:0] core_io_dmem_resp_bits_data; // @[top.scala 21:26]
  wire  core__GEN_451; // @[top.scala 21:26]
  wire  core__GEN_331; // @[top.scala 21:26]
  wire  core__GEN_337; // @[top.scala 21:26]
  wire  core__GEN_113; // @[top.scala 21:26]
  wire  core__GEN_111; // @[top.scala 21:26]
  wire  core__GEN_415; // @[top.scala 21:26]
  wire  core__GEN_436; // @[top.scala 21:26]
  wire  core__GEN_140; // @[top.scala 21:26]
  wire  core__GEN_71; // @[top.scala 21:26]
  wire  core__GEN_324; // @[top.scala 21:26]
  wire  core__GEN_219; // @[top.scala 21:26]
  wire  core__GEN_168; // @[top.scala 21:26]
  wire  core__GEN_98; // @[top.scala 21:26]
  wire  core__GEN_1; // @[top.scala 21:26]
  wire  core__GEN_352; // @[top.scala 21:26]
  wire  core__GEN_423; // @[top.scala 21:26]
  wire  core__GEN_44; // @[top.scala 21:26]
  wire  core__GEN_125; // @[top.scala 21:26]
  wire  core__GEN_267; // @[top.scala 21:26]
  wire  core__GEN_126; // @[top.scala 21:26]
  wire  core__GEN_430; // @[top.scala 21:26]
  wire  core__GEN_153; // @[top.scala 21:26]
  wire  core__GEN_225; // @[top.scala 21:26]
  wire  core__GEN_119; // @[top.scala 21:26]
  wire  core__GEN_88; // @[top.scala 21:26]
  wire  core__GEN_59; // @[top.scala 21:26]
  wire  core__GEN_252; // @[top.scala 21:26]
  wire  core__GEN_151; // @[top.scala 21:26]
  wire  core__GEN_147; // @[top.scala 21:26]
  wire  core__GEN_310; // @[top.scala 21:26]
  wire  core__GEN_351; // @[top.scala 21:26]
  wire  core__GEN_210; // @[top.scala 21:26]
  wire  core__GEN_246; // @[top.scala 21:26]
  wire  core__GEN_104; // @[top.scala 21:26]
  wire  core__GEN_409; // @[top.scala 21:26]
  wire  core__GEN_65; // @[top.scala 21:26]
  wire  core__GEN_253; // @[top.scala 21:26]
  wire  core__GEN_132; // @[top.scala 21:26]
  wire  core__GEN_318; // @[top.scala 21:26]
  wire  core__GEN_316; // @[top.scala 21:26]
  wire  core__GEN_92; // @[top.scala 21:26]
  wire  core__GEN_345; // @[top.scala 21:26]
  wire  core__GEN_231; // @[top.scala 21:26]
  wire  core__GEN_417; // @[top.scala 21:26]
  wire  core__GEN_244; // @[top.scala 21:26]
  wire  core__GEN_50; // @[top.scala 21:26]
  wire  core__GEN_238; // @[top.scala 21:26]
  wire  core__GEN_330; // @[top.scala 21:26]
  wire  core__GEN_86; // @[top.scala 21:26]
  wire  core__GEN_339; // @[top.scala 21:26]
  wire  core__GEN_101; // @[top.scala 21:26]
  wire  core__GEN_325; // @[top.scala 21:26]
  wire  core__GEN_240; // @[top.scala 21:26]
  wire  core__GEN_234; // @[top.scala 21:26]
  wire  core__GEN_120; // @[top.scala 21:26]
  wire  core__GEN_169; // @[top.scala 21:26]
  wire  core__GEN_129; // @[top.scala 21:26]
  wire  core__GEN_433; // @[top.scala 21:26]
  wire  core__GEN_333; // @[top.scala 21:26]
  wire  core__GEN_302; // @[top.scala 21:26]
  wire  core__GEN_313; // @[top.scala 21:26]
  wire  core__GEN_228; // @[top.scala 21:26]
  wire  core__GEN_197; // @[top.scala 21:26]
  wire  core__GEN_91; // @[top.scala 21:26]
  wire  core__GEN_411; // @[top.scala 21:26]
  wire  core__GEN_11; // @[top.scala 21:26]
  wire  core__GEN_401; // @[top.scala 21:26]
  wire  core__GEN_47; // @[top.scala 21:26]
  wire  core__GEN_296; // @[top.scala 21:26]
  wire  core__GEN_304; // @[top.scala 21:26]
  wire  core__GEN_294; // @[top.scala 21:26]
  wire  core__GEN_74; // @[top.scala 21:26]
  wire  core__GEN_213; // @[top.scala 21:26]
  wire  core__GEN_303; // @[top.scala 21:26]
  wire  core__GEN_107; // @[top.scala 21:26]
  wire  core__GEN_32; // @[top.scala 21:26]
  wire  core__GEN_0; // @[top.scala 21:26]
  wire  core__GEN_402; // @[top.scala 21:26]
  wire  core__GEN_412; // @[top.scala 21:26]
  wire  core__GEN_68; // @[top.scala 21:26]
  wire  core__GEN_135; // @[top.scala 21:26]
  wire  core__GEN_424; // @[top.scala 21:26]
  wire  core__GEN_175; // @[top.scala 21:26]
  wire  core__GEN_319; // @[top.scala 21:26]
  wire  core__GEN_288; // @[top.scala 21:26]
  wire  core__GEN_56; // @[top.scala 21:26]
  wire  core__GEN_26; // @[top.scala 21:26]
  wire  core__GEN_418; // @[top.scala 21:26]
  wire  core__GEN_122; // @[top.scala 21:26]
  wire  core__GEN_387; // @[top.scala 21:26]
  wire  core__GEN_53; // @[top.scala 21:26]
  wire  core__GEN_141; // @[top.scala 21:26]
  wire  core__GEN_327; // @[top.scala 21:26]
  wire  core__GEN_72; // @[top.scala 21:26]
  wire  core__GEN_395; // @[top.scala 21:26]
  wire  core__GEN_249; // @[top.scala 21:26]
  wire  core__GEN_114; // @[top.scala 21:26]
  wire  core__GEN_312; // @[top.scala 21:26]
  wire  core__GEN_203; // @[top.scala 21:26]
  wire  core__GEN_75; // @[top.scala 21:26]
  wire  core__GEN_85; // @[top.scala 21:26]
  wire  core__GEN_20; // @[top.scala 21:26]
  wire  core__GEN_178; // @[top.scala 21:26]
  wire  core__GEN_15; // @[top.scala 21:26]
  wire  core__GEN_157; // @[top.scala 21:26]
  wire  core__GEN_462; // @[top.scala 21:26]
  wire  core__GEN_69; // @[top.scala 21:26]
  wire  core__GEN_216; // @[top.scala 21:26]
  wire  core__GEN_206; // @[top.scala 21:26]
  wire  core__GEN_375; // @[top.scala 21:26]
  wire  core__GEN_151_0; // @[top.scala 21:26]
  wire  core__GEN_420; // @[top.scala 21:26]
  wire  core__GEN_123; // @[top.scala 21:26]
  wire  core__GEN_315; // @[top.scala 21:26]
  wire  core__GEN_284; // @[top.scala 21:26]
  wire  core__GEN_179; // @[top.scala 21:26]
  wire  core__GEN_33; // @[top.scala 21:26]
  wire  core__GEN_222; // @[top.scala 21:26]
  wire  core__GEN_377; // @[top.scala 21:26]
  wire  core__GEN_191; // @[top.scala 21:26]
  wire  core__GEN_290; // @[top.scala 21:26]
  wire  core__GEN_404; // @[top.scala 21:26]
  wire  core__GEN_390; // @[top.scala 21:26]
  wire  core__GEN_56_0; // @[top.scala 21:26]
  wire  core__GEN_305; // @[top.scala 21:26]
  wire  core__GEN_299; // @[top.scala 21:26]
  wire  core__GEN_185; // @[top.scala 21:26]
  wire  core__GEN_307; // @[top.scala 21:26]
  wire  core__GEN_297; // @[top.scala 21:26]
  wire  core__GEN_398; // @[top.scala 21:26]
  wire  core__GEN_406; // @[top.scala 21:26]
  wire  core__GEN_41; // @[top.scala 21:26]
  wire  core__GEN_321; // @[top.scala 21:26]
  wire  core__GEN_270; // @[top.scala 21:26]
  wire  core__GEN_95; // @[top.scala 21:26]
  wire  core__GEN_45; // @[top.scala 21:26]
  wire  core__GEN_414; // @[top.scala 21:26]
  wire  core__GEN_383; // @[top.scala 21:26]
  wire  core__GEN_369; // @[top.scala 21:26]
  wire  core__GEN_35; // @[top.scala 21:26]
  wire  core__GEN_29; // @[top.scala 21:26]
  wire  core__GEN_278; // @[top.scala 21:26]
  wire  core__GEN_117; // @[top.scala 21:26]
  wire  core__GEN_396; // @[top.scala 21:26]
  wire  core__GEN_172; // @[top.scala 21:26]
  wire  core__GEN_276; // @[top.scala 21:26]
  wire  core__GEN_291; // @[top.scala 21:26]
  wire  core__GEN_365; // @[top.scala 21:26]
  wire  core__GEN_359; // @[top.scala 21:26]
  wire  core__GEN_258; // @[top.scala 21:26]
  wire  core__GEN_372; // @[top.scala 21:26]
  wire  core__GEN_38; // @[top.scala 21:26]
  wire  core__GEN_252_0; // @[top.scala 21:26]
  wire  core__GEN_167; // @[top.scala 21:26]
  wire  core__GEN_166; // @[top.scala 21:26]
  wire  core__GEN_285; // @[top.scala 21:26]
  wire  core__GEN_42; // @[top.scala 21:26]
  wire  core__GEN_350; // @[top.scala 21:26]
  wire  core__GEN_106; // @[top.scala 21:26]
  wire  core__GEN_384; // @[top.scala 21:26]
  wire  core__GEN_18; // @[top.scala 21:26]
  wire  core__GEN_378; // @[top.scala 21:26]
  wire  core__GEN_393; // @[top.scala 21:26]
  wire  core__GEN_273; // @[top.scala 21:26]
  wire  core__GEN_293; // @[top.scala 21:26]
  wire  core__GEN_456; // @[top.scala 21:26]
  wire  core__GEN_371; // @[top.scala 21:26]
  wire  core__GEN_80; // @[top.scala 21:26]
  wire  core__GEN_351_0; // @[top.scala 21:26]
  wire  core__GEN_251; // @[top.scala 21:26]
  wire  core__GEN_209; // @[top.scala 21:26]
  wire  core__GEN_139; // @[top.scala 21:26]
  wire  core__GEN_145; // @[top.scala 21:26]
  wire  core__GEN_450; // @[top.scala 21:26]
  wire  core__GEN_308; // @[top.scala 21:26]
  wire  core__GEN_173; // @[top.scala 21:26]
  wire  core__GEN_53_0; // @[top.scala 21:26]
  wire  core__GEN_357; // @[top.scala 21:26]
  wire  core__GEN_200; // @[top.scala 21:26]
  wire  core__GEN_386; // @[top.scala 21:26]
  wire  core__GEN_272; // @[top.scala 21:26]
  wire  core__GEN_160; // @[top.scala 21:26]
  wire  core__GEN_91_0; // @[top.scala 21:26]
  wire  core__GEN_279; // @[top.scala 21:26]
  wire  core__GEN_194; // @[top.scala 21:26]
  wire  core__GEN_188; // @[top.scala 21:26]
  wire  core__GEN_133; // @[top.scala 21:26]
  wire  core__GEN_392; // @[top.scala 21:26]
  wire  core__GEN_23; // @[top.scala 21:26]
  wire  core__GEN_407; // @[top.scala 21:26]
  wire  core__GEN_287; // @[top.scala 21:26]
  wire  core__GEN_266; // @[top.scala 21:26]
  wire  core__GEN_399; // @[top.scala 21:26]
  wire  core__GEN_264; // @[top.scala 21:26]
  wire  core__GEN_300; // @[top.scala 21:26]
  wire  core__GEN_374; // @[top.scala 21:26]
  wire  core__GEN_233; // @[top.scala 21:26]
  wire  core__GEN_127; // @[top.scala 21:26]
  wire  core__GEN_269; // @[top.scala 21:26]
  wire  core__GEN_432; // @[top.scala 21:26]
  wire  core__GEN_381; // @[top.scala 21:26]
  wire  core__GEN_260; // @[top.scala 21:26]
  wire  core__GEN_161; // @[top.scala 21:26]
  wire  core__GEN_155; // @[top.scala 21:26]
  wire  core__GEN_339_0; // @[top.scala 21:26]
  wire  core__GEN_368; // @[top.scala 21:26]
  wire  core__GEN_254; // @[top.scala 21:26]
  wire  core__GEN_281; // @[top.scala 21:26]
  wire  core__GEN_73; // @[top.scala 21:26]
  wire  core__GEN_261; // @[top.scala 21:26]
  wire  core__GEN_353; // @[top.scala 21:26]
  wire  core__GEN_332; // @[top.scala 21:26]
  wire  core__GEN_88_0; // @[top.scala 21:26]
  wire  core__GEN_176; // @[top.scala 21:26]
  wire  core__GEN_16; // @[top.scala 21:26]
  wire  core__GEN_380; // @[top.scala 21:26]
  wire  core__GEN_360; // @[top.scala 21:26]
  wire  core__GEN_389; // @[top.scala 21:26]
  wire  core__GEN_163; // @[top.scala 21:26]
  wire  core__GEN_246_0; // @[top.scala 21:26]
  wire  core__GEN_438; // @[top.scala 21:26]
  wire  core__GEN_94; // @[top.scala 21:26]
  wire  core__GEN_282; // @[top.scala 21:26]
  wire  core__GEN_347; // @[top.scala 21:26]
  wire  core__GEN_109; // @[top.scala 21:26]
  wire  core__GEN_182; // @[top.scala 21:26]
  wire  core__GEN_345_0; // @[top.scala 21:26]
  wire  core__GEN_121; // @[top.scala 21:26]
  wire  core__GEN_240_0; // @[top.scala 21:26]
  wire  core__GEN_9; // @[top.scala 21:26]
  wire  core__GEN_148; // @[top.scala 21:26]
  wire  core__GEN_154; // @[top.scala 21:26]
  wire  core__GEN_444; // @[top.scala 21:26]
  wire  core__GEN_149; // @[top.scala 21:26]
  wire  core__GEN_267_0; // @[top.scala 21:26]
  wire  core__GEN_459; // @[top.scala 21:26]
  wire  core__GEN_453; // @[top.scala 21:26]
  wire  core__GEN_248; // @[top.scala 21:26]
  wire  core__GEN_366; // @[top.scala 21:26]
  wire  core__GEN_7; // @[top.scala 21:26]
  wire  core__GEN_142; // @[top.scala 21:26]
  wire  core__GEN_275; // @[top.scala 21:26]
  wire  core__GEN_140_0; // @[top.scala 21:26]
  wire  core__GEN_324_0; // @[top.scala 21:26]
  wire  core__GEN_100; // @[top.scala 21:26]
  wire  core__GEN_333_0; // @[top.scala 21:26]
  wire  core__GEN_362; // @[top.scala 21:26]
  wire  core__GEN_413; // @[top.scala 21:26]
  wire  core__GEN_342; // @[top.scala 21:26]
  wire  core__GEN_405; // @[top.scala 21:26]
  wire  core__GEN_420_0; // @[top.scala 21:26]
  wire  core__GEN_306; // @[top.scala 21:26]
  wire  core__GEN_76; // @[top.scala 21:26]
  wire  core__GEN_164; // @[top.scala 21:26]
  wire  core__GEN_109_0; // @[top.scala 21:26]
  wire  core__GEN_103; // @[top.scala 21:26]
  wire  core__GEN_3; // @[top.scala 21:26]
  wire  core__GEN_242; // @[top.scala 21:26]
  wire  core__GEN_136; // @[top.scala 21:26]
  wire  core__GEN_426; // @[top.scala 21:26]
  wire  core__GEN_137; // @[top.scala 21:26]
  wire  core__GEN_441; // @[top.scala 21:26]
  wire  core__GEN_341; // @[top.scala 21:26]
  wire  core__GEN_94_0; // @[top.scala 21:26]
  wire  core__GEN_348; // @[top.scala 21:26]
  wire  core__GEN_263; // @[top.scala 21:26]
  wire  core__GEN_257; // @[top.scala 21:26]
  wire  core__GEN_122_0; // @[top.scala 21:26]
  wire  core__GEN_143; // @[top.scala 21:26]
  wire  core__GEN_255; // @[top.scala 21:26]
  wire  core__GEN_82; // @[top.scala 21:26]
  wire  core__GEN_170; // @[top.scala 21:26]
  wire  core__GEN_356; // @[top.scala 21:26]
  wire  core__GEN_221; // @[top.scala 21:26]
  wire  core__GEN_215; // @[top.scala 21:26]
  wire  core__GEN_115; // @[top.scala 21:26]
  wire  core__GEN_146; // @[top.scala 21:26]
  wire  core__GEN_363; // @[top.scala 21:26]
  wire  core__GEN_320; // @[top.scala 21:26]
  wire  core__GEN_314; // @[top.scala 21:26]
  wire  core__GEN_329; // @[top.scala 21:26]
  wire  core__GEN_321_0; // @[top.scala 21:26]
  wire  core__GEN_327_0; // @[top.scala 21:26]
  wire  core__GEN_103_0; // @[top.scala 21:26]
  wire  core__GEN_97; // @[top.scala 21:26]
  wire  core__GEN_236; // @[top.scala 21:26]
  wire  core__GEN_354; // @[top.scala 21:26]
  wire  core__GEN_234_0; // @[top.scala 21:26]
  wire  core__GEN_130; // @[top.scala 21:26]
  wire  core__GEN_61; // @[top.scala 21:26]
  wire  core__GEN_55; // @[top.scala 21:26]
  wire  core__GEN_249_0; // @[top.scala 21:26]
  wire  core__GEN_335; // @[top.scala 21:26]
  wire  core__GEN_243; // @[top.scala 21:26]
  wire  core__GEN_447; // @[top.scala 21:26]
  wire  core__GEN_158; // @[top.scala 21:26]
  wire  core__GEN_330_0; // @[top.scala 21:26]
  wire  core__GEN_422; // @[top.scala 21:26]
  wire  core__GEN_245; // @[top.scala 21:26]
  wire  core__GEN_37; // @[top.scala 21:26]
  wire  core__GEN_125_0; // @[top.scala 21:26]
  wire  core__GEN_429; // @[top.scala 21:26]
  wire  core__GEN_70; // @[top.scala 21:26]
  wire  core__GEN_64; // @[top.scala 21:26]
  wire  core__GEN_344; // @[top.scala 21:26]
  wire  core__GEN_338; // @[top.scala 21:26]
  wire  core__GEN_293_0; // @[top.scala 21:26]
  wire  core__GEN_87; // @[top.scala 21:26]
  wire  core__GEN_416; // @[top.scala 21:26]
  wire  core__GEN_406_0; // @[top.scala 21:26]
  wire  core__GEN_58; // @[top.scala 21:26]
  wire  core__GEN_414_0; // @[top.scala 21:26]
  wire  core__GEN_309; // @[top.scala 21:26]
  wire  core__GEN_85_0; // @[top.scala 21:26]
  wire  core__GEN_299_0; // @[top.scala 21:26]
  wire  core__GEN_336; // @[top.scala 21:26]
  wire  core__GEN_408; // @[top.scala 21:26]
  wire  core__GEN_112; // @[top.scala 21:26]
  wire  core__GEN_43; // @[top.scala 21:26]
  wire  core__GEN_150; // @[top.scala 21:26]
  wire  core__GEN_131; // @[top.scala 21:26]
  wire  core__GEN_435; // @[top.scala 21:26]
  wire  core__GEN_230; // @[top.scala 21:26]
  wire  core__GEN_97_0; // @[top.scala 21:26]
  wire  core__GEN_124; // @[top.scala 21:26]
  wire  core__GEN_239; // @[top.scala 21:26]
  wire  core__GEN_118; // @[top.scala 21:26]
  wire  core__GEN_392_0; // @[top.scala 21:26]
  wire  core__GEN_398_0; // @[top.scala 21:26]
  wire  core__GEN_423_0; // @[top.scala 21:26]
  wire  core__GEN_237; // @[top.scala 21:26]
  wire  core__GEN_152; // @[top.scala 21:26]
  wire  core__GEN_307_0; // @[top.scala 21:26]
  wire  core__GEN_146_0; // @[top.scala 21:26]
  wire  core__GEN_315_0; // @[top.scala 21:26]
  wire  core__GEN_79; // @[top.scala 21:26]
  wire  core__GEN_224; // @[top.scala 21:26]
  wire  core__GEN_110; // @[top.scala 21:26]
  wire  core__GEN_119_0; // @[top.scala 21:26]
  wire  core__GEN_323; // @[top.scala 21:26]
  wire  core__GEN_317; // @[top.scala 21:26]
  wire  core__GEN_79_0; // @[top.scala 21:26]
  wire  core__GEN_218; // @[top.scala 21:26]
  wire  core__GEN_208; // @[top.scala 21:26]
  wire  core__GEN_1_1; // @[top.scala 21:26]
  wire  core__GEN_196; // @[top.scala 21:26]
  wire  core__GEN_90; // @[top.scala 21:26]
  wire  core__GEN_31; // @[top.scala 21:26]
  wire  core__GEN_400; // @[top.scala 21:26]
  wire  core__GEN_113_0; // @[top.scala 21:26]
  wire  core__GEN_162; // @[top.scala 21:26]
  wire  core__GEN_212; // @[top.scala 21:26]
  wire  core__GEN_302_0; // @[top.scala 21:26]
  wire  core__GEN_181; // @[top.scala 21:26]
  wire  core__GEN_106_0; // @[top.scala 21:26]
  wire  core__GEN_227; // @[top.scala 21:26]
  wire  core__GEN_71_0; // @[top.scala 21:26]
  wire  core__GEN_380_0; // @[top.scala 21:26]
  wire  core__GEN_425; // @[top.scala 21:26]
  wire  core__GEN_280; // @[top.scala 21:26]
  wire  core__GEN_46; // @[top.scala 21:26]
  wire  core__GEN_174; // @[top.scala 21:26]
  wire  core__GEN_134; // @[top.scala 21:26]
  wire  core__GEN_289; // @[top.scala 21:26]
  wire  core__GEN_318_0; // @[top.scala 21:26]
  wire  core__GEN_287_0; // @[top.scala 21:26]
  wire  core__GEN_202; // @[top.scala 21:26]
  wire  core__GEN_419; // @[top.scala 21:26]
  wire  core__GEN_388; // @[top.scala 21:26]
  wire  core__GEN_410; // @[top.scala 21:26]
  wire  core__GEN_386_0; // @[top.scala 21:26]
  wire  core__GEN_52; // @[top.scala 21:26]
  wire  core__GEN_311; // @[top.scala 21:26]
  wire  core__GEN_301; // @[top.scala 21:26]
  wire  core__GEN_295; // @[top.scala 21:26]
  wire  core__GEN_67; // @[top.scala 21:26]
  wire  core__GEN_281_0; // @[top.scala 21:26]
  wire  core__GEN_312_0; // @[top.scala 21:26]
  wire  core__GEN_25; // @[top.scala 21:26]
  wire  core__GEN_409_0; // @[top.scala 21:26]
  wire  core__GEN_417_0; // @[top.scala 21:26]
  wire  core__GEN_411_0; // @[top.scala 21:26]
  wire  core__GEN_326; // @[top.scala 21:26]
  wire  core__GEN_55_0; // @[top.scala 21:26]
  wire  core__GEN_100_0; // @[top.scala 21:26]
  wire  core__GEN_394; // @[top.scala 21:26]
  wire  core__GEN_168_0; // @[top.scala 21:26]
  wire  core__GEN_128; // @[top.scala 21:26]
  wire  core__GEN_401_0; // @[top.scala 21:26]
  wire  core__GEN_44_0; // @[top.scala 21:26]
  wire  core__GEN_376; // @[top.scala 21:26]
  wire  core__GEN_74_0; // @[top.scala 21:26]
  wire  core__GEN_374_0; // @[top.scala 21:26]
  wire  core__GEN_40; // @[top.scala 21:26]
  wire  core__GEN_368_0; // @[top.scala 21:26]
  wire  core__GEN_34; // @[top.scala 21:26]
  wire  core__GEN_383_0; // @[top.scala 21:26]
  wire  core__GEN_49; // @[top.scala 21:26]
  wire  core__GEN_263_0; // @[top.scala 21:26]
  wire  core__GEN_177; // @[top.scala 21:26]
  wire  core__GEN_171; // @[top.scala 21:26]
  wire  core__GEN_446; // @[top.scala 21:26]
  wire  core__GEN_102; // @[top.scala 21:26]
  wire  core__GEN_290_0; // @[top.scala 21:26]
  wire  core__GEN_190; // @[top.scala 21:26]
  wire  core__GEN_83; // @[top.scala 21:26]
  wire  core__GEN_205; // @[top.scala 21:26]
  wire  core__GEN_135_0; // @[top.scala 21:26]
  wire  core__GEN_389_0; // @[top.scala 21:26]
  wire  core__GEN_93; // @[top.scala 21:26]
  wire  core__GEN_254_0; // @[top.scala 21:26]
  wire  core__GEN_298; // @[top.scala 21:26]
  wire  core__GEN_163_0; // @[top.scala 21:26]
  wire  core__GEN_21; // @[top.scala 21:26]
  wire  core__GEN_461; // @[top.scala 21:26]
  wire  core__GEN_362_0; // @[top.scala 21:26]
  wire  core__GEN_14; // @[top.scala 21:26]
  wire  core__GEN_116; // @[top.scala 21:26]
  wire  core__GEN_156; // @[top.scala 21:26]
  wire  core__GEN_150_0; // @[top.scala 21:26]
  wire  core__GEN_283; // @[top.scala 21:26]
  wire  core__GEN_184; // @[top.scala 21:26]
  wire  core__GEN_178_0; // @[top.scala 21:26]
  wire  core__GEN_68_0; // @[top.scala 21:26]
  wire  core__GEN_296_0; // @[top.scala 21:26]
  wire  core__GEN_382; // @[top.scala 21:26]
  wire  core__GEN_397; // @[top.scala 21:26]
  wire  core__GEN_277; // @[top.scala 21:26]
  wire  core__GEN_395_0; // @[top.scala 21:26]
  wire  core__GEN_304_0; // @[top.scala 21:26]
  wire  core__GEN_199; // @[top.scala 21:26]
  wire  core__GEN_403; // @[top.scala 21:26]
  wire  core__GEN_262; // @[top.scala 21:26]
  wire  core__GEN_28; // @[top.scala 21:26]
  wire  core__GEN_275_0; // @[top.scala 21:26]
  wire  core__GEN_269_0; // @[top.scala 21:26]
  wire  core__GEN_361; // @[top.scala 21:26]
  wire  core__GEN_96; // @[top.scala 21:26]
  wire  core__GEN_278_0; // @[top.scala 21:26]
  wire  core__GEN_193; // @[top.scala 21:26]
  wire  core__GEN_379; // @[top.scala 21:26]
  wire  core__GEN_244_0; // @[top.scala 21:26]
  wire  core__GEN_138; // @[top.scala 21:26]
  wire  core__GEN_271; // @[top.scala 21:26]
  wire  core__GEN_251_0; // @[top.scala 21:26]
  wire  core__GEN_151_1; // @[top.scala 21:26]
  wire  core__GEN_166_0; // @[top.scala 21:26]
  wire  core__GEN_455; // @[top.scala 21:26]
  wire  core__GEN_370; // @[top.scala 21:26]
  wire  core__GEN_364; // @[top.scala 21:26]
  wire  core__GEN_259; // @[top.scala 21:26]
  wire  core__GEN_377_0; // @[top.scala 21:26]
  wire  core__GEN_153_0; // @[top.scala 21:26]
  wire  core__GEN_292; // @[top.scala 21:26]
  wire  core__GEN_84; // @[top.scala 21:26]
  wire  core__GEN_78; // @[top.scala 21:26]
  wire  core__GEN_272_0; // @[top.scala 21:26]
  wire  core__GEN_47_0; // @[top.scala 21:26]
  wire  core__GEN_335_0; // @[top.scala 21:26]
  wire  core__GEN_41_0; // @[top.scala 21:26]
  wire  core__GEN_385; // @[top.scala 21:26]
  wire  core__GEN_250; // @[top.scala 21:26]
  wire  core__GEN_434; // @[top.scala 21:26]
  wire  core__GEN_257_0; // @[top.scala 21:26]
  wire  core__GEN_343; // @[top.scala 21:26]
  wire  core__GEN_443; // @[top.scala 21:26]
  wire  core__GEN_105; // @[top.scala 21:26]
  wire  core__GEN_99; // @[top.scala 21:26]
  wire  core__GEN_358; // @[top.scala 21:26]
  wire  core__GEN_356_0; // @[top.scala 21:26]
  wire  core__GEN_350_0; // @[top.scala 21:26]
  wire  core__GEN_132_0; // @[top.scala 21:26]
  wire  core__GEN_22; // @[top.scala 21:26]
  wire  core__GEN_144; // @[top.scala 21:26]
  wire  core__GEN_265; // @[top.scala 21:26]
  wire  core__GEN_17; // @[top.scala 21:26]
  wire  core__GEN_159; // @[top.scala 21:26]
  wire  core__GEN_428; // @[top.scala 21:26]
  wire  core__GEN_449; // @[top.scala 21:26]
  wire  core__GEN_90_0; // @[top.scala 21:26]
  wire  core__GEN_172_0; // @[top.scala 21:26]
  wire  core__GEN_187; // @[top.scala 21:26]
  wire  core__GEN_117_0; // @[top.scala 21:26]
  wire  core__GEN_236_0; // @[top.scala 21:26]
  wire  core__GEN_371_0; // @[top.scala 21:26]
  wire  core__GEN_391; // @[top.scala 21:26]
  wire  core__GEN_165; // @[top.scala 21:26]
  wire  core__GEN_286; // @[top.scala 21:26]
  wire  core__GEN_145_0; // @[top.scala 21:26]
  wire  core__GEN_284_0; // @[top.scala 21:26]
  wire  core__GEN_232; // @[top.scala 21:26]
  wire  core__GEN_147_0; // @[top.scala 21:26]
  wire  core__GEN_416_0; // @[top.scala 21:26]
  wire  core__GEN_274; // @[top.scala 21:26]
  wire  core__GEN_260_0; // @[top.scala 21:26]
  wire  core__GEN_175_0; // @[top.scala 21:26]
  wire  core__GEN_105_0; // @[top.scala 21:26]
  wire  core__GEN_169_0; // @[top.scala 21:26]
  wire  core__GEN_338_0; // @[top.scala 21:26]
  wire  core__GEN_247; // @[top.scala 21:26]
  wire  core__GEN_133_0; // @[top.scala 21:26]
  wire  core__GEN_141_0; // @[top.scala 21:26]
  wire  core__GEN_160_0; // @[top.scala 21:26]
  wire  core__GEN_346; // @[top.scala 21:26]
  wire  core__GEN_99_0; // @[top.scala 21:26]
  wire  core__GEN_344_0; // @[top.scala 21:26]
  wire  core__GEN_373; // @[top.scala 21:26]
  wire  core__GEN_424_0; // @[top.scala 21:26]
  wire  core__GEN_239_0; // @[top.scala 21:26]
  wire  core__GEN_353_0; // @[top.scala 21:26]
  wire  core__GEN_268; // @[top.scala 21:26]
  wire  core__GEN_127_0; // @[top.scala 21:26]
  wire  core__GEN_8; // @[top.scala 21:26]
  wire  core__GEN_266_0; // @[top.scala 21:26]
  wire  core__GEN_331_0; // @[top.scala 21:26]
  wire  core__GEN_452; // @[top.scala 21:26]
  wire  core__GEN_93_0; // @[top.scala 21:26]
  wire  core__GEN_87_0; // @[top.scala 21:26]
  wire  core__GEN_367; // @[top.scala 21:26]
  wire  core__GEN_226; // @[top.scala 21:26]
  wire  core__GEN_120_0; // @[top.scala 21:26]
  wire  core__GEN_365_0; // @[top.scala 21:26]
  wire  core__GEN_6; // @[top.scala 21:26]
  wire  core__GEN_410_0; // @[top.scala 21:26]
  wire  core__GEN_253_0; // @[top.scala 21:26]
  wire  core__GEN_152_0; // @[top.scala 21:26]
  wire  core__GEN_325_0; // @[top.scala 21:26]
  wire  core__GEN_148_0; // @[top.scala 21:26]
  wire  core__GEN_437; // @[top.scala 21:26]
  wire  core__GEN_352_0; // @[top.scala 21:26]
  wire  core__GEN_332_0; // @[top.scala 21:26]
  wire  core__GEN_108; // @[top.scala 21:26]
  wire  core__GEN_126_0; // @[top.scala 21:26]
  wire  core__GEN_245_0; // @[top.scala 21:26]
  wire  core__GEN_359_0; // @[top.scala 21:26]
  wire  core__GEN_431; // @[top.scala 21:26]
  wire  core__GEN_72_0; // @[top.scala 21:26]
  wire  core__GEN_66; // @[top.scala 21:26]
  wire  core__GEN_154_0; // @[top.scala 21:26]
  wire  core__GEN_458; // @[top.scala 21:26]
  wire  core__GEN_317_0; // @[top.scala 21:26]
  wire  core__GEN_326_0; // @[top.scala 21:26]
  wire  core__GEN_241; // @[top.scala 21:26]
  wire  core__GEN_341_0; // @[top.scala 21:26]
  wire  core__GEN_402_0; // @[top.scala 21:26]
  wire  core__GEN_1_2; // @[top.scala 21:26]
  wire  core__GEN_48; // @[top.scala 21:26]
  wire  core__GEN_394_0; // @[top.scala 21:26]
  wire  core__GEN_60; // @[top.scala 21:26]
  wire  core__GEN_248_0; // @[top.scala 21:26]
  wire  core__GEN_75_0; // @[top.scala 21:26]
  wire  core__GEN_349; // @[top.scala 21:26]
  wire  core__GEN_214; // @[top.scala 21:26]
  wire  core__GEN_347_0; // @[top.scala 21:26]
  wire  core__GEN_412_0; // @[top.scala 21:26]
  wire  core__GEN_92_0; // @[top.scala 21:26]
  wire  core__GEN_102_0; // @[top.scala 21:26]
  wire  core__GEN_256; // @[top.scala 21:26]
  wire  core__GEN_121_0; // @[top.scala 21:26]
  wire  core__GEN_425_0; // @[top.scala 21:26]
  wire  core__GEN_305_0; // @[top.scala 21:26]
  wire  core__GEN_419_0; // @[top.scala 21:26]
  wire  core__GEN_81; // @[top.scala 21:26]
  wire  core__GEN_320_0; // @[top.scala 21:26]
  wire  core__GEN_108_0; // @[top.scala 21:26]
  wire  core__GEN_114_0; // @[top.scala 21:26]
  wire  core__GEN_123_0; // @[top.scala 21:26]
  wire  core__GEN_413_0; // @[top.scala 21:26]
  wire  core__GEN_54; // @[top.scala 21:26]
  wire  core__GEN_136_0; // @[top.scala 21:26]
  wire  core__GEN_142_0; // @[top.scala 21:26]
  wire  core__GEN_440; // @[top.scala 21:26]
  wire  core__GEN_295_0; // @[top.scala 21:26]
  wire  core__GEN_340; // @[top.scala 21:26]
  wire  core__GEN_355; // @[top.scala 21:26]
  wire  core__GEN_235; // @[top.scala 21:26]
  wire  core__GEN_129_0; // @[top.scala 21:26]
  wire  core__GEN_404_0; // @[top.scala 21:26]
  wire  core__GEN_403_0; // @[top.scala 21:26]
  wire  core__GEN_313_0; // @[top.scala 21:26]
  wire  core__GEN_242_0; // @[top.scala 21:26]
  wire  core__GEN_69_0; // @[top.scala 21:26]
  wire  core__GEN_157_0; // @[top.scala 21:26]
  wire  core__GEN_220; // @[top.scala 21:26]
  wire  core__GEN_229; // @[top.scala 21:26]
  wire  core__GEN_115_0; // @[top.scala 21:26]
  wire  core__GEN_15_0; // @[top.scala 21:26]
  wire  core__GEN_334; // @[top.scala 21:26]
  wire  core__GEN_328; // @[top.scala 21:26]
  wire  core__GEN_96_0; // @[top.scala 21:26]
  wire  core__GEN_86_0; // @[top.scala 21:26]
  wire  core__GEN_36; // @[top.scala 21:26]
  wire  core__GEN_405_0; // @[top.scala 21:26]
  wire  core__GEN_415_0; // @[top.scala 21:26]
  wire  core__GEN_164_0; // @[top.scala 21:26]
  wire  core__GEN_124_0; // @[top.scala 21:26]
  wire  core__GEN_322; // @[top.scala 21:26]
  wire  core__GEN_308_0; // @[top.scala 21:26]
  wire  core__GEN_337_0; // @[top.scala 21:26]
  wire  core__GEN_223; // @[top.scala 21:26]
  wire  core__GEN_217; // @[top.scala 21:26]
  wire  core__GEN_192; // @[top.scala 21:26]
  wire  core__GEN_390_0; // @[top.scala 21:26]
  wire  core__GEN_42_0; // @[top.scala 21:26]
  wire  core__GEN_149_0; // @[top.scala 21:26]
  wire  core__GEN_291_0; // @[top.scala 21:26]
  wire  core__GEN_139_0; // @[top.scala 21:26]
  wire  core__GEN_329_0; // @[top.scala 21:26]
  wire  core__GEN_292_0; // @[top.scala 21:26]
  wire  core__GEN_298_0; // @[top.scala 21:26]
  wire  core__GEN_207; // @[top.scala 21:26]
  wire  core__GEN_399_0; // @[top.scala 21:26]
  wire  core__GEN_421; // @[top.scala 21:26]
  wire  core__GEN_63; // @[top.scala 21:26]
  wire  core__GEN_391_0; // @[top.scala 21:26]
  wire  core__GEN_316_0; // @[top.scala 21:26]
  wire  core__GEN_306_0; // @[top.scala 21:26]
  wire  core__GEN_314_0; // @[top.scala 21:26]
  wire  core__GEN_21_0; // @[top.scala 21:26]
  wire  core__GEN_323_0; // @[top.scala 21:26]
  wire  core__GEN_384_0; // @[top.scala 21:26]
  wire  core__GEN_118_0; // @[top.scala 21:26]
  wire  core__GEN_376_0; // @[top.scala 21:26]
  wire  core__GEN_422_0; // @[top.scala 21:26]
  wire  core__GEN_277_0; // @[top.scala 21:26]
  wire  core__GEN_57; // @[top.scala 21:26]
  wire  core__GEN_130_0; // @[top.scala 21:26]
  wire  core__GEN_46_0; // @[top.scala 21:26]
  wire  core__GEN_111_0; // @[top.scala 21:26]
  wire  core__GEN_78_0; // @[top.scala 21:26]
  wire  core__GEN_238_0; // @[top.scala 21:26]
  wire  core__GEN_407_0; // @[top.scala 21:26]
  wire  core__GEN_179_0; // @[top.scala 21:26]
  wire  core__GEN_397_0; // @[top.scala 21:26]
  wire  core__GEN_173_0; // @[top.scala 21:26]
  wire  core__GEN_70_0; // @[top.scala 21:26]
  wire  core__GEN_379_0; // @[top.scala 21:26]
  wire  core__GEN_82_0; // @[top.scala 21:26]
  wire  core__GEN_373_0; // @[top.scala 21:26]
  wire  core__GEN_45_0; // @[top.scala 21:26]
  wire  core__GEN_54_0; // @[top.scala 21:26]
  wire  core__GEN_201; // @[top.scala 21:26]
  wire  core__GEN_195; // @[top.scala 21:26]
  wire  core__GEN_364_0; // @[top.scala 21:26]
  wire  core__GEN_259_0; // @[top.scala 21:26]
  wire  core__GEN_167_0; // @[top.scala 21:26]
  wire  core__GEN_309_0; // @[top.scala 21:26]
  wire  core__GEN_43_0; // @[top.scala 21:26]
  wire  core__GEN_372_0; // @[top.scala 21:26]
  wire  core__GEN_19; // @[top.scala 21:26]
  wire  core__GEN_161_0; // @[top.scala 21:26]
  wire  core__GEN_51; // @[top.scala 21:26]
  wire  core__GEN_265_0; // @[top.scala 21:26]
  wire  core__GEN_294_0; // @[top.scala 21:26]
  wire  core__GEN_180; // @[top.scala 21:26]
  wire  core__GEN_189; // @[top.scala 21:26]
  wire  core__GEN_211; // @[top.scala 21:26]
  wire  core__GEN_301_0; // @[top.scala 21:26]
  wire  core__GEN_393_0; // @[top.scala 21:26]
  wire  core__GEN_387_0; // @[top.scala 21:26]
  wire  core__GEN_39; // @[top.scala 21:26]
  wire  core__GEN_146_1; // @[top.scala 21:26]
  wire  core__GEN_288_0; // @[top.scala 21:26]
  wire  core__GEN_310_0; // @[top.scala 21:26]
  wire  core__GEN_300_0; // @[top.scala 21:26]
  wire  core__GEN_286_0; // @[top.scala 21:26]
  wire  core__GEN_400_0; // @[top.scala 21:26]
  wire  core__GEN_319_0; // @[top.scala 21:26]
  wire  core__GEN_107_0; // @[top.scala 21:26]
  wire  core__GEN_174_0; // @[top.scala 21:26]
  wire  core__GEN_89; // @[top.scala 21:26]
  wire  core__GEN_358_0; // @[top.scala 21:26]
  wire  core__GEN_30; // @[top.scala 21:26]
  wire  core__GEN_24; // @[top.scala 21:26]
  wire  core__GEN_408_0; // @[top.scala 21:26]
  wire  core__GEN_418_0; // @[top.scala 21:26]
  wire  core__GEN_273_0; // @[top.scala 21:26]
  wire  core__GEN_5_0; // @[top.scala 21:26]
  wire  core__GEN_112_0; // @[top.scala 21:26]
  wire  core__GEN_385_0; // @[top.scala 21:26]
  wire  core__GEN_457; // @[top.scala 21:26]
  wire  core__GEN_311_0; // @[top.scala 21:26]
  wire  core__GEN_280_0; // @[top.scala 21:26]
  wire  core__GEN_366_0; // @[top.scala 21:26]
  wire  core__GEN_360_0; // @[top.scala 21:26]
  wire  core__GEN_354_0; // @[top.scala 21:26]
  wire  core__GEN_143_0; // @[top.scala 21:26]
  wire  core__GEN_367_0; // @[top.scala 21:26]
  wire  core__GEN_33_0; // @[top.scala 21:26]
  wire  core__GEN_247_0; // @[top.scala 21:26]
  wire  core__GEN_276_0; // @[top.scala 21:26]
  wire  core__GEN_348_0; // @[top.scala 21:26]
  wire  core__GEN_274_0; // @[top.scala 21:26]
  wire  core__GEN_460; // @[top.scala 21:26]
  wire  core__GEN_101_0; // @[top.scala 21:26]
  wire  core__GEN_375_0; // @[top.scala 21:26]
  wire  core__GEN_283_0; // @[top.scala 21:26]
  wire  core__GEN_27; // @[top.scala 21:26]
  wire  core__GEN_13; // @[top.scala 21:26]
  wire  core__GEN_388_0; // @[top.scala 21:26]
  wire  core__GEN_382_0; // @[top.scala 21:26]
  wire  core__GEN_268_0; // @[top.scala 21:26]
  wire  core__GEN_297_0; // @[top.scala 21:26]
  wire  core__GEN_89_0; // @[top.scala 21:26]
  wire  core__GEN_176_0; // @[top.scala 21:26]
  wire  core__GEN_177_0; // @[top.scala 21:26]
  wire  core__GEN_346_0; // @[top.scala 21:26]
  wire  core__GEN_64_0; // @[top.scala 21:26]
  wire  core__GEN_340_0; // @[top.scala 21:26]
  wire  core__GEN_255_0; // @[top.scala 21:26]
  wire  core__GEN_204; // @[top.scala 21:26]
  wire  core__GEN_134_0; // @[top.scala 21:26]
  wire  core__GEN_149_1; // @[top.scala 21:26]
  wire  core__GEN_439; // @[top.scala 21:26]
  wire  core__GEN_80_0; // @[top.scala 21:26]
  wire  core__GEN_262_0; // @[top.scala 21:26]
  wire  core__GEN_303_0; // @[top.scala 21:26]
  wire  core__GEN_162_0; // @[top.scala 21:26]
  wire  core__GEN_17_0; // @[top.scala 21:26]
  wire  core__GEN_198; // @[top.scala 21:26]
  wire  core__GEN_361_0; // @[top.scala 21:26]
  wire  core__GEN_381_0; // @[top.scala 21:26]
  wire  core__GEN_261_0; // @[top.scala 21:26]
  wire  core__GEN_155_0; // @[top.scala 21:26]
  wire  core__GEN_156_0; // @[top.scala 21:26]
  wire  core__GEN_170_0; // @[top.scala 21:26]
  wire  core__GEN_95_0; // @[top.scala 21:26]
  wire  core__GEN_183; // @[top.scala 21:26]
  wire  core__GEN_369_0; // @[top.scala 21:26]
  wire  core__GEN_73_0; // @[top.scala 21:26]
  wire  core__GEN_128_0; // @[top.scala 21:26]
  wire  core__GEN_241_0; // @[top.scala 21:26]
  wire  core__GEN_282_0; // @[top.scala 21:26]
  wire  core__GEN_396_0; // @[top.scala 21:26]
  wire  core__GEN_445; // @[top.scala 21:26]
  wire  core__GEN_289_0; // @[top.scala 21:26]
  wire  core__GEN_378_0; // @[top.scala 21:26]
  wire  core__GEN_186; // @[top.scala 21:26]
  wire  core__GEN_131_0; // @[top.scala 21:26]
  wire  core__GEN_152_1; // @[top.scala 21:26]
  wire  core__GEN_421_0; // @[top.scala 21:26]
  wire  core__GEN_427; // @[top.scala 21:26]
  wire  core__GEN_62; // @[top.scala 21:26]
  wire  core__GEN_285_0; // @[top.scala 21:26]
  wire  core__GEN_336_0; // @[top.scala 21:26]
  wire  core__GEN_144_0; // @[top.scala 21:26]
  wire  core__GEN_150_1; // @[top.scala 21:26]
  wire  core__GEN_454; // @[top.scala 21:26]
  wire  core__GEN_363_0; // @[top.scala 21:26]
  wire  core__GEN_243_0; // @[top.scala 21:26]
  wire  core__GEN_258_0; // @[top.scala 21:26]
  wire  core__GEN_138_0; // @[top.scala 21:26]
  wire  core__GEN_256_0; // @[top.scala 21:26]
  wire  core__GEN_171_0; // @[top.scala 21:26]
  wire  core__GEN_357_0; // @[top.scala 21:26]
  wire  core__GEN_165_0; // @[top.scala 21:26]
  wire  core__GEN_110_0; // @[top.scala 21:26]
  wire  core__GEN_40_0; // @[top.scala 21:26]
  wire  core__GEN_264_0; // @[top.scala 21:26]
  wire  core__GEN_5_1; // @[top.scala 21:26]
  wire  core__GEN_158_0; // @[top.scala 21:26]
  wire  core__GEN_16_0; // @[top.scala 21:26]
  wire  core__GEN_271_0; // @[top.scala 21:26]
  wire  core__GEN_342_0; // @[top.scala 21:26]
  wire  core__GEN_322_0; // @[top.scala 21:26]
  wire  core__GEN_98_0; // @[top.scala 21:26]
  wire  core__GEN_237_0; // @[top.scala 21:26]
  wire  core__GEN_334_0; // @[top.scala 21:26]
  wire  core__GEN_116_0; // @[top.scala 21:26]
  wire  core__GEN_235_0; // @[top.scala 21:26]
  wire  core__GEN_349_0; // @[top.scala 21:26]
  wire  core__GEN_147_1; // @[top.scala 21:26]
  wire  core__GEN_448; // @[top.scala 21:26]
  wire  core__GEN_442; // @[top.scala 21:26]
  wire  core__GEN_83_0; // @[top.scala 21:26]
  wire  core__GEN_343_0; // @[top.scala 21:26]
  wire  core__GEN_355_0; // @[top.scala 21:26]
  wire  core__GEN_137_0; // @[top.scala 21:26]
  wire  core__GEN_370_0; // @[top.scala 21:26]
  wire  core__GEN_250_0; // @[top.scala 21:26]
  wire  core__GEN_77; // @[top.scala 21:26]
  wire  core__GEN_270_0; // @[top.scala 21:26]
  wire  core__GEN_279_0; // @[top.scala 21:26]
  wire  core__GEN_159_0; // @[top.scala 21:26]
  wire  core__GEN_463; // @[top.scala 21:26]
  wire  core__GEN_328_0; // @[top.scala 21:26]
  wire  core__GEN_104_0; // @[top.scala 21:26]
  wire  memory_metaReset; // @[top.scala 24:28]
  wire  memory_clock; // @[top.scala 24:28]
  wire  memory_io_core_ports_0_req_valid; // @[top.scala 24:28]
  wire [31:0] memory_io_core_ports_0_req_bits_addr; // @[top.scala 24:28]
  wire [31:0] memory_io_core_ports_0_req_bits_data; // @[top.scala 24:28]
  wire  memory_io_core_ports_0_req_bits_fcn; // @[top.scala 24:28]
  wire [2:0] memory_io_core_ports_0_req_bits_typ; // @[top.scala 24:28]
  wire  memory_io_core_ports_0_resp_valid; // @[top.scala 24:28]
  wire [31:0] memory_io_core_ports_0_resp_bits_data; // @[top.scala 24:28]
  wire  memory__GEN_4_0; // @[top.scala 24:28]
  wire  memory__GEN_1_1; // @[top.scala 24:28]
  wire  memory__GEN_0_1; // @[top.scala 24:28]
  wire  memory__GEN_3_1; // @[top.scala 24:28]
  wire  memory__GEN_5_0; // @[top.scala 24:28]
  wire  memory__GEN_2_0; // @[top.scala 24:28]
  wire  profilePin = core__GEN_1;
  wire  profilePin_0 = core__GEN_5_0;
  wire  profilePin_1 = core__GEN_8;
  wire  profilePin_2 = core__GEN_9;
  wire  profilePin_3 = core__GEN_13;
  wire  profilePin_4 = core__GEN_14;
  wire  profilePin_5 = core__GEN_15;
  wire  profilePin_6 = core__GEN_16_0;
  wire  profilePin_7 = core__GEN_17;
  wire  profilePin_8 = core__GEN_18;
  wire [9:0] _GEN_803 = {profilePin,profilePin_0,profilePin_1,profilePin_2,profilePin_3,profilePin_4,profilePin_5,profilePin_6,profilePin_7,profilePin_8};
  wire  profilePin_9 = core__GEN_19;
  wire  profilePin_10 = core__GEN_20;
  wire  profilePin_11 = core__GEN_21_0;
  wire  profilePin_12 = core__GEN_22;
  wire  profilePin_13 = core__GEN_23;
  wire  profilePin_14 = core__GEN_24;
  wire  profilePin_15 = core__GEN_25;
  wire  profilePin_16 = core__GEN_26;
  wire  profilePin_17 = core__GEN_27;
  wire [18:0] _GEN_812 = {_GEN_803,profilePin_9,profilePin_10,profilePin_11,profilePin_12,profilePin_13,profilePin_14,profilePin_15,profilePin_16,profilePin_17};
  wire  profilePin_18 = core__GEN_28;
  wire  profilePin_19 = core__GEN_29;
  wire  profilePin_20 = core__GEN_30;
  wire  profilePin_21 = core__GEN_31;
  wire  profilePin_22 = core__GEN_32;
  wire  profilePin_23 = core__GEN_33_0;
  wire  profilePin_24 = core__GEN_34;
  wire  profilePin_25 = core__GEN_35;
  wire  profilePin_26 = core__GEN_36;
  wire [27:0] _GEN_821 = {_GEN_812,profilePin_18,profilePin_19,profilePin_20,profilePin_21,profilePin_22,profilePin_23,profilePin_24,profilePin_25,profilePin_26};
  wire  profilePin_27 = core__GEN_37;
  wire  profilePin_28 = core__GEN_38;
  wire  profilePin_29 = core__GEN_39;
  wire  profilePin_30 = core__GEN_40;
  wire  profilePin_31 = core__GEN_41;
  wire  profilePin_32 = core__GEN_42_0;
  wire  profilePin_33 = core__GEN_43;
  wire  profilePin_34 = core__GEN_44;
  wire  profilePin_35 = core__GEN_45_0;
  wire [36:0] _GEN_830 = {_GEN_821,profilePin_27,profilePin_28,profilePin_29,profilePin_30,profilePin_31,profilePin_32,profilePin_33,profilePin_34,profilePin_35};
  wire  profilePin_36 = core__GEN_46;
  wire  profilePin_37 = core__GEN_47;
  wire  profilePin_38 = core__GEN_48;
  wire  profilePin_39 = core__GEN_49;
  wire  profilePin_40 = core__GEN_50;
  wire  profilePin_41 = core__GEN_51;
  wire  profilePin_42 = core__GEN_52;
  wire  profilePin_43 = core__GEN_53;
  wire  profilePin_44 = core__GEN_54;
  wire [45:0] _GEN_839 = {_GEN_830,profilePin_36,profilePin_37,profilePin_38,profilePin_39,profilePin_40,profilePin_41,profilePin_42,profilePin_43,profilePin_44};
  wire  profilePin_45 = core__GEN_55;
  wire  profilePin_46 = core__GEN_56_0;
  wire  profilePin_47 = core__GEN_57;
  wire  profilePin_48 = core__GEN_58;
  wire  profilePin_49 = core__GEN_59;
  wire  profilePin_50 = core__GEN_60;
  wire  profilePin_51 = core__GEN_61;
  wire  profilePin_52 = core__GEN_62;
  wire  profilePin_53 = core__GEN_63;
  wire [54:0] _GEN_848 = {_GEN_839,profilePin_45,profilePin_46,profilePin_47,profilePin_48,profilePin_49,profilePin_50,profilePin_51,profilePin_52,profilePin_53};
  wire  profilePin_54 = core__GEN_64;
  wire  profilePin_55 = core__GEN_65;
  wire  profilePin_56 = core__GEN_66;
  wire  profilePin_57 = core__GEN_67;
  wire  profilePin_58 = core__GEN_68;
  wire  profilePin_59 = core__GEN_69_0;
  wire  profilePin_60 = core__GEN_70;
  wire  profilePin_61 = core__GEN_71;
  wire  profilePin_62 = core__GEN_72_0;
  wire [63:0] _GEN_857 = {_GEN_848,profilePin_54,profilePin_55,profilePin_56,profilePin_57,profilePin_58,profilePin_59,profilePin_60,profilePin_61,profilePin_62};
  wire  profilePin_63 = core__GEN_73;
  wire  profilePin_64 = core__GEN_74;
  wire  profilePin_65 = core__GEN_75_0;
  wire  profilePin_66 = core__GEN_76;
  wire  profilePin_67 = core__GEN_77;
  wire  profilePin_68 = core__GEN_78;
  wire  profilePin_69 = core__GEN_79_0;
  wire  profilePin_70 = core__GEN_80_0;
  wire  profilePin_71 = core__GEN_81;
  wire [72:0] _GEN_866 = {_GEN_857,profilePin_63,profilePin_64,profilePin_65,profilePin_66,profilePin_67,profilePin_68,profilePin_69,profilePin_70,profilePin_71};
  wire  profilePin_72 = core__GEN_82;
  wire  profilePin_73 = core__GEN_83_0;
  wire  profilePin_74 = core__GEN_84;
  wire  profilePin_75 = core__GEN_85_0;
  wire  profilePin_76 = core__GEN_86;
  wire  profilePin_77 = core__GEN_87_0;
  wire  profilePin_78 = core__GEN_88_0;
  wire  profilePin_79 = core__GEN_89_0;
  wire  profilePin_80 = core__GEN_90_0;
  wire [81:0] _GEN_875 = {_GEN_866,profilePin_72,profilePin_73,profilePin_74,profilePin_75,profilePin_76,profilePin_77,profilePin_78,profilePin_79,profilePin_80};
  wire  profilePin_81 = core__GEN_91_0;
  wire  profilePin_82 = core__GEN_92;
  wire  profilePin_83 = core__GEN_93_0;
  wire  profilePin_84 = core__GEN_94;
  wire  profilePin_85 = core__GEN_95_0;
  wire  profilePin_86 = core__GEN_96;
  wire  profilePin_87 = core__GEN_97;
  wire  profilePin_88 = core__GEN_98_0;
  wire  profilePin_89 = core__GEN_99;
  wire [90:0] _GEN_884 = {_GEN_875,profilePin_81,profilePin_82,profilePin_83,profilePin_84,profilePin_85,profilePin_86,profilePin_87,profilePin_88,profilePin_89};
  wire  profilePin_90 = core__GEN_100;
  wire  profilePin_91 = core__GEN_101_0;
  wire  profilePin_92 = core__GEN_102;
  wire  profilePin_93 = core__GEN_103_0;
  wire  profilePin_94 = core__GEN_104_0;
  wire  profilePin_95 = core__GEN_105;
  wire  profilePin_96 = core__GEN_106;
  wire  profilePin_97 = core__GEN_107_0;
  wire  profilePin_98 = core__GEN_108;
  wire [99:0] _GEN_893 = {_GEN_884,profilePin_90,profilePin_91,profilePin_92,profilePin_93,profilePin_94,profilePin_95,profilePin_96,profilePin_97,profilePin_98};
  wire  profilePin_99 = core__GEN_109;
  wire  profilePin_100 = core__GEN_110;
  wire  profilePin_101 = core__GEN_111;
  wire  profilePin_102 = core__GEN_112_0;
  wire  profilePin_103 = core__GEN_113_0;
  wire  profilePin_104 = core__GEN_114;
  wire  profilePin_105 = core__GEN_115_0;
  wire  profilePin_106 = core__GEN_116;
  wire  profilePin_107 = core__GEN_117;
  wire [108:0] _GEN_902 = {_GEN_893,profilePin_99,profilePin_100,profilePin_101,profilePin_102,profilePin_103,profilePin_104,profilePin_105,profilePin_106,profilePin_107};
  wire  profilePin_108 = core__GEN_118_0;
  wire  profilePin_109 = core__GEN_119_0;
  wire  profilePin_110 = core__GEN_120;
  wire  profilePin_111 = core__GEN_121_0;
  wire  profilePin_112 = core__GEN_122_0;
  wire  profilePin_113 = core__GEN_123;
  wire  profilePin_114 = core__GEN_124_0;
  wire  profilePin_115 = core__GEN_125_0;
  wire  profilePin_116 = core__GEN_126;
  wire [117:0] _GEN_911 = {_GEN_902,profilePin_108,profilePin_109,profilePin_110,profilePin_111,profilePin_112,profilePin_113,profilePin_114,profilePin_115,profilePin_116};
  wire  profilePin_117 = core__GEN_127_0;
  wire  profilePin_118 = core__GEN_128;
  wire  profilePin_119 = core__GEN_129;
  wire  profilePin_120 = core__GEN_130_0;
  wire  profilePin_121 = core__GEN_131;
  wire  profilePin_122 = core__GEN_132;
  wire  profilePin_123 = core__GEN_133_0;
  wire  profilePin_124 = core__GEN_134;
  wire  profilePin_125 = core__GEN_135;
  wire [126:0] _GEN_920 = {_GEN_911,profilePin_117,profilePin_118,profilePin_119,profilePin_120,profilePin_121,profilePin_122,profilePin_123,profilePin_124,profilePin_125};
  wire  profilePin_126 = core__GEN_136_0;
  wire  profilePin_127 = core__GEN_137;
  wire  profilePin_128 = core__GEN_138_0;
  wire  profilePin_129 = core__GEN_139_0;
  wire  profilePin_130 = core__GEN_140_0;
  wire  profilePin_131 = core__GEN_141;
  wire  profilePin_132 = core__GEN_142_0;
  wire  profilePin_133 = core__GEN_143;
  wire  profilePin_134 = core__GEN_144_0;
  wire [135:0] _GEN_929 = {_GEN_920,profilePin_126,profilePin_127,profilePin_128,profilePin_129,profilePin_130,profilePin_131,profilePin_132,profilePin_133,profilePin_134};
  wire  profilePin_135 = core__GEN_145_0;
  wire  profilePin_136 = core__GEN_146_0;
  wire  profilePin_137 = core__GEN_147;
  wire  profilePin_138 = core__GEN_148_0;
  wire  profilePin_139 = core__GEN_149;
  wire  profilePin_140 = core__GEN_150_1;
  wire  profilePin_141 = core__GEN_151_1;
  wire  profilePin_142 = core__GEN_152;
  wire  profilePin_143 = core__GEN_153;
  wire [144:0] _GEN_938 = {_GEN_929,profilePin_135,profilePin_136,profilePin_137,profilePin_138,profilePin_139,profilePin_140,profilePin_141,profilePin_142,profilePin_143};
  wire  profilePin_144 = core__GEN_154_0;
  wire  profilePin_145 = core__GEN_155;
  wire  profilePin_146 = core__GEN_156_0;
  wire  profilePin_147 = core__GEN_157_0;
  wire  profilePin_148 = core__GEN_158;
  wire  profilePin_149 = core__GEN_159_0;
  wire  profilePin_150 = core__GEN_160_0;
  wire  profilePin_151 = core__GEN_161;
  wire  profilePin_152 = core__GEN_162_0;
  wire [153:0] _GEN_947 = {_GEN_938,profilePin_144,profilePin_145,profilePin_146,profilePin_147,profilePin_148,profilePin_149,profilePin_150,profilePin_151,profilePin_152};
  wire  profilePin_153 = core__GEN_163_0;
  wire  profilePin_154 = core__GEN_164;
  wire  profilePin_155 = core__GEN_165_0;
  wire  profilePin_156 = core__GEN_166_0;
  wire  profilePin_157 = core__GEN_167;
  wire  profilePin_158 = core__GEN_168;
  wire  profilePin_159 = core__GEN_169_0;
  wire  profilePin_160 = core__GEN_170;
  wire  profilePin_161 = core__GEN_171_0;
  wire [162:0] _GEN_956 = {_GEN_947,profilePin_153,profilePin_154,profilePin_155,profilePin_156,profilePin_157,profilePin_158,profilePin_159,profilePin_160,profilePin_161};
  wire  profilePin_162 = core__GEN_172_0;
  wire  profilePin_163 = core__GEN_173;
  wire  profilePin_164 = core__GEN_174_0;
  wire  profilePin_165 = core__GEN_175_0;
  wire  profilePin_166 = core__GEN_176;
  wire  profilePin_167 = core__GEN_177_0;
  wire  profilePin_168 = core__GEN_178_0;
  wire  profilePin_169 = core__GEN_179;
  wire  profilePin_170 = core__GEN_180;
  wire [171:0] _GEN_965 = {_GEN_956,profilePin_162,profilePin_163,profilePin_164,profilePin_165,profilePin_166,profilePin_167,profilePin_168,profilePin_169,profilePin_170};
  wire  profilePin_171 = core__GEN_181;
  wire  profilePin_172 = core__GEN_182;
  wire  profilePin_173 = core__GEN_183;
  wire  profilePin_174 = core__GEN_184;
  wire  profilePin_175 = core__GEN_185;
  wire  profilePin_176 = core__GEN_186;
  wire  profilePin_177 = core__GEN_187;
  wire  profilePin_178 = core__GEN_188;
  wire  profilePin_179 = core__GEN_189;
  wire [180:0] _GEN_974 = {_GEN_965,profilePin_171,profilePin_172,profilePin_173,profilePin_174,profilePin_175,profilePin_176,profilePin_177,profilePin_178,profilePin_179};
  wire  profilePin_180 = core__GEN_190;
  wire  profilePin_181 = core__GEN_191;
  wire  profilePin_182 = core__GEN_192;
  wire  profilePin_183 = core__GEN_193;
  wire  profilePin_184 = core__GEN_194;
  wire  profilePin_185 = core__GEN_195;
  wire  profilePin_186 = core__GEN_196;
  wire  profilePin_187 = core__GEN_197;
  wire  profilePin_188 = core__GEN_198;
  wire [189:0] _GEN_983 = {_GEN_974,profilePin_180,profilePin_181,profilePin_182,profilePin_183,profilePin_184,profilePin_185,profilePin_186,profilePin_187,profilePin_188};
  wire  profilePin_189 = core__GEN_199;
  wire  profilePin_190 = core__GEN_200;
  wire  profilePin_191 = core__GEN_201;
  wire  profilePin_192 = core__GEN_202;
  wire  profilePin_193 = core__GEN_203;
  wire  profilePin_194 = core__GEN_204;
  wire  profilePin_195 = core__GEN_205;
  wire  profilePin_196 = core__GEN_206;
  wire  profilePin_197 = core__GEN_207;
  wire [198:0] _GEN_992 = {_GEN_983,profilePin_189,profilePin_190,profilePin_191,profilePin_192,profilePin_193,profilePin_194,profilePin_195,profilePin_196,profilePin_197};
  wire  profilePin_198 = core__GEN_208;
  wire  profilePin_199 = core__GEN_209;
  wire  profilePin_200 = core__GEN_210;
  wire  profilePin_201 = core__GEN_211;
  wire  profilePin_202 = core__GEN_212;
  wire  profilePin_203 = core__GEN_213;
  wire  profilePin_204 = core__GEN_214;
  wire  profilePin_205 = core__GEN_215;
  wire  profilePin_206 = core__GEN_216;
  wire [207:0] _GEN_1001 = {_GEN_992,profilePin_198,profilePin_199,profilePin_200,profilePin_201,profilePin_202,profilePin_203,profilePin_204,profilePin_205,profilePin_206};
  wire  profilePin_207 = core__GEN_217;
  wire  profilePin_208 = core__GEN_218;
  wire  profilePin_209 = core__GEN_219;
  wire  profilePin_210 = core__GEN_220;
  wire  profilePin_211 = core__GEN_221;
  wire  profilePin_212 = core__GEN_222;
  wire  profilePin_213 = core__GEN_223;
  wire  profilePin_214 = core__GEN_224;
  wire  profilePin_215 = core__GEN_225;
  wire [216:0] _GEN_1010 = {_GEN_1001,profilePin_207,profilePin_208,profilePin_209,profilePin_210,profilePin_211,profilePin_212,profilePin_213,profilePin_214,profilePin_215};
  wire  profilePin_216 = core__GEN_226;
  wire  profilePin_217 = core__GEN_227;
  wire  profilePin_218 = core__GEN_228;
  wire  profilePin_219 = core__GEN_229;
  wire  profilePin_220 = core__GEN_230;
  wire  profilePin_221 = core__GEN_231;
  wire  profilePin_222 = core__GEN_232;
  wire  profilePin_223 = core__GEN_233;
  wire  profilePin_224 = core__GEN_234;
  wire [225:0] _GEN_1019 = {_GEN_1010,profilePin_216,profilePin_217,profilePin_218,profilePin_219,profilePin_220,profilePin_221,profilePin_222,profilePin_223,profilePin_224};
  wire  profilePin_225 = core__GEN_235;
  wire  profilePin_226 = core__GEN_236;
  wire  profilePin_227 = core__GEN_237_0;
  wire  profilePin_228 = core__GEN_238_0;
  wire  profilePin_229 = core__GEN_239;
  wire  profilePin_230 = core__GEN_240;
  wire  profilePin_231 = core__GEN_241;
  wire  profilePin_232 = core__GEN_242;
  wire  profilePin_233 = core__GEN_243_0;
  wire [234:0] _GEN_1028 = {_GEN_1019,profilePin_225,profilePin_226,profilePin_227,profilePin_228,profilePin_229,profilePin_230,profilePin_231,profilePin_232,profilePin_233};
  wire  profilePin_234 = core__GEN_244_0;
  wire  profilePin_235 = core__GEN_245;
  wire  profilePin_236 = core__GEN_246;
  wire  profilePin_237 = core__GEN_247;
  wire  profilePin_238 = core__GEN_248;
  wire  profilePin_239 = core__GEN_249;
  wire  profilePin_240 = core__GEN_250;
  wire  profilePin_241 = core__GEN_251;
  wire  profilePin_242 = core__GEN_252;
  wire [243:0] _GEN_1037 = {_GEN_1028,profilePin_234,profilePin_235,profilePin_236,profilePin_237,profilePin_238,profilePin_239,profilePin_240,profilePin_241,profilePin_242};
  wire  profilePin_243 = core__GEN_253_0;
  wire  profilePin_244 = core__GEN_254;
  wire  profilePin_245 = core__GEN_255_0;
  wire  profilePin_246 = core__GEN_256;
  wire  profilePin_247 = core__GEN_257;
  wire  profilePin_248 = core__GEN_258_0;
  wire  profilePin_249 = core__GEN_259;
  wire  profilePin_250 = core__GEN_260;
  wire  profilePin_251 = core__GEN_261_0;
  wire [252:0] _GEN_1046 = {_GEN_1037,profilePin_243,profilePin_244,profilePin_245,profilePin_246,profilePin_247,profilePin_248,profilePin_249,profilePin_250,profilePin_251};
  wire  profilePin_252 = core__GEN_262;
  wire  profilePin_253 = core__GEN_263;
  wire  profilePin_254 = core__GEN_264_0;
  wire  profilePin_255 = core__GEN_265;
  wire  profilePin_256 = core__GEN_266;
  wire  profilePin_257 = core__GEN_267;
  wire  profilePin_258 = core__GEN_268;
  wire  profilePin_259 = core__GEN_269;
  wire  profilePin_260 = core__GEN_270_0;
  wire [261:0] _GEN_1055 = {_GEN_1046,profilePin_252,profilePin_253,profilePin_254,profilePin_255,profilePin_256,profilePin_257,profilePin_258,profilePin_259,profilePin_260};
  wire  profilePin_261 = core__GEN_271;
  wire  profilePin_262 = core__GEN_272;
  wire  profilePin_263 = core__GEN_273_0;
  wire  profilePin_264 = core__GEN_274;
  wire  profilePin_265 = core__GEN_275;
  wire  profilePin_266 = core__GEN_276_0;
  wire  profilePin_267 = core__GEN_277;
  wire  profilePin_268 = core__GEN_278;
  wire  profilePin_269 = core__GEN_279_0;
  wire [270:0] _GEN_1064 = {_GEN_1055,profilePin_261,profilePin_262,profilePin_263,profilePin_264,profilePin_265,profilePin_266,profilePin_267,profilePin_268,profilePin_269};
  wire  profilePin_270 = core__GEN_280;
  wire  profilePin_271 = core__GEN_281;
  wire  profilePin_272 = core__GEN_282_0;
  wire  profilePin_273 = core__GEN_283;
  wire  profilePin_274 = core__GEN_284;
  wire  profilePin_275 = core__GEN_285_0;
  wire  profilePin_276 = core__GEN_286;
  wire  profilePin_277 = core__GEN_287;
  wire  profilePin_278 = core__GEN_288_0;
  wire [279:0] _GEN_1073 = {_GEN_1064,profilePin_270,profilePin_271,profilePin_272,profilePin_273,profilePin_274,profilePin_275,profilePin_276,profilePin_277,profilePin_278};
  wire  profilePin_279 = core__GEN_289;
  wire  profilePin_280 = core__GEN_290;
  wire  profilePin_281 = core__GEN_291_0;
  wire  profilePin_282 = core__GEN_292;
  wire  profilePin_283 = core__GEN_293;
  wire  profilePin_284 = core__GEN_294_0;
  wire  profilePin_285 = core__GEN_295;
  wire  profilePin_286 = core__GEN_296;
  wire  profilePin_287 = core__GEN_297_0;
  wire [288:0] _GEN_1082 = {_GEN_1073,profilePin_279,profilePin_280,profilePin_281,profilePin_282,profilePin_283,profilePin_284,profilePin_285,profilePin_286,profilePin_287};
  wire  profilePin_288 = core__GEN_298;
  wire  profilePin_289 = core__GEN_299;
  wire  profilePin_290 = core__GEN_300_0;
  wire  profilePin_291 = core__GEN_301;
  wire  profilePin_292 = core__GEN_302;
  wire  profilePin_293 = core__GEN_303_0;
  wire  profilePin_294 = core__GEN_304_0;
  wire  profilePin_295 = core__GEN_305;
  wire  profilePin_296 = core__GEN_306_0;
  wire [297:0] _GEN_1091 = {_GEN_1082,profilePin_288,profilePin_289,profilePin_290,profilePin_291,profilePin_292,profilePin_293,profilePin_294,profilePin_295,profilePin_296};
  wire  profilePin_297 = core__GEN_307_0;
  wire  profilePin_298 = core__GEN_308;
  wire  profilePin_299 = core__GEN_309_0;
  wire  profilePin_300 = core__GEN_310_0;
  wire  profilePin_301 = core__GEN_311;
  wire  profilePin_302 = core__GEN_312;
  wire  profilePin_303 = core__GEN_313_0;
  wire  profilePin_304 = core__GEN_314;
  wire  profilePin_305 = core__GEN_315;
  wire [306:0] _GEN_1100 = {_GEN_1091,profilePin_297,profilePin_298,profilePin_299,profilePin_300,profilePin_301,profilePin_302,profilePin_303,profilePin_304,profilePin_305};
  wire  profilePin_306 = core__GEN_316_0;
  wire  profilePin_307 = core__GEN_317;
  wire  profilePin_308 = core__GEN_318;
  wire  profilePin_309 = core__GEN_319_0;
  wire  profilePin_310 = core__GEN_320;
  wire  profilePin_311 = core__GEN_321;
  wire  profilePin_312 = core__GEN_322;
  wire  profilePin_313 = core__GEN_323;
  wire  profilePin_314 = core__GEN_324;
  wire [315:0] _GEN_1109 = {_GEN_1100,profilePin_306,profilePin_307,profilePin_308,profilePin_309,profilePin_310,profilePin_311,profilePin_312,profilePin_313,profilePin_314};
  wire  profilePin_315 = core__GEN_325_0;
  wire  profilePin_316 = core__GEN_326;
  wire  profilePin_317 = core__GEN_327;
  wire  profilePin_318 = core__GEN_328;
  wire  profilePin_319 = core__GEN_329;
  wire  profilePin_320 = core__GEN_330;
  wire  profilePin_321 = core__GEN_331_0;
  wire  profilePin_322 = core__GEN_332;
  wire  profilePin_323 = core__GEN_333;
  wire [324:0] _GEN_1118 = {_GEN_1109,profilePin_315,profilePin_316,profilePin_317,profilePin_318,profilePin_319,profilePin_320,profilePin_321,profilePin_322,profilePin_323};
  wire  profilePin_324 = core__GEN_334;
  wire  profilePin_325 = core__GEN_335;
  wire  profilePin_326 = core__GEN_336_0;
  wire  profilePin_327 = core__GEN_337_0;
  wire  profilePin_328 = core__GEN_338;
  wire  profilePin_329 = core__GEN_339;
  wire  profilePin_330 = core__GEN_340;
  wire  profilePin_331 = core__GEN_341;
  wire  profilePin_332 = core__GEN_342_0;
  wire [333:0] _GEN_1127 = {_GEN_1118,profilePin_324,profilePin_325,profilePin_326,profilePin_327,profilePin_328,profilePin_329,profilePin_330,profilePin_331,profilePin_332};
  wire  profilePin_333 = core__GEN_343;
  wire  profilePin_334 = core__GEN_344;
  wire  profilePin_335 = core__GEN_345;
  wire  profilePin_336 = core__GEN_346;
  wire  profilePin_337 = core__GEN_347;
  wire  profilePin_338 = core__GEN_348_0;
  wire  profilePin_339 = core__GEN_349;
  wire  profilePin_340 = core__GEN_350;
  wire  profilePin_341 = core__GEN_351;
  wire [342:0] _GEN_1136 = {_GEN_1127,profilePin_333,profilePin_334,profilePin_335,profilePin_336,profilePin_337,profilePin_338,profilePin_339,profilePin_340,profilePin_341};
  wire  profilePin_342 = core__GEN_352_0;
  wire  profilePin_343 = core__GEN_353;
  wire  profilePin_344 = core__GEN_354_0;
  wire  profilePin_345 = core__GEN_355;
  wire  profilePin_346 = core__GEN_356;
  wire  profilePin_347 = core__GEN_357_0;
  wire  profilePin_348 = core__GEN_358;
  wire  profilePin_349 = core__GEN_359;
  wire  profilePin_350 = core__GEN_360_0;
  wire [351:0] _GEN_1145 = {_GEN_1136,profilePin_342,profilePin_343,profilePin_344,profilePin_345,profilePin_346,profilePin_347,profilePin_348,profilePin_349,profilePin_350};
  wire  profilePin_351 = core__GEN_361;
  wire  profilePin_352 = core__GEN_362;
  wire  profilePin_353 = core__GEN_363_0;
  wire  profilePin_354 = core__GEN_364;
  wire  profilePin_355 = core__GEN_365;
  wire  profilePin_356 = core__GEN_366_0;
  wire  profilePin_357 = core__GEN_367;
  wire  profilePin_358 = core__GEN_368;
  wire  profilePin_359 = core__GEN_369_0;
  wire [360:0] _GEN_1154 = {_GEN_1145,profilePin_351,profilePin_352,profilePin_353,profilePin_354,profilePin_355,profilePin_356,profilePin_357,profilePin_358,profilePin_359};
  wire  profilePin_360 = core__GEN_370;
  wire  profilePin_361 = core__GEN_371;
  wire  profilePin_362 = core__GEN_372_0;
  wire  profilePin_363 = core__GEN_373;
  wire  profilePin_364 = core__GEN_374;
  wire  profilePin_365 = core__GEN_375_0;
  wire  profilePin_366 = core__GEN_376;
  wire  profilePin_367 = core__GEN_377;
  wire  profilePin_368 = core__GEN_378_0;
  wire [369:0] _GEN_1163 = {_GEN_1154,profilePin_360,profilePin_361,profilePin_362,profilePin_363,profilePin_364,profilePin_365,profilePin_366,profilePin_367,profilePin_368};
  wire  profilePin_369 = core__GEN_379;
  wire  profilePin_370 = core__GEN_380;
  wire  profilePin_371 = core__GEN_381_0;
  wire  profilePin_372 = core__GEN_382;
  wire  profilePin_373 = core__GEN_383;
  wire  profilePin_374 = core__GEN_384_0;
  wire  profilePin_375 = core__GEN_385;
  wire  profilePin_376 = core__GEN_386;
  wire  profilePin_377 = core__GEN_387_0;
  wire [378:0] _GEN_1172 = {_GEN_1163,profilePin_369,profilePin_370,profilePin_371,profilePin_372,profilePin_373,profilePin_374,profilePin_375,profilePin_376,profilePin_377};
  wire  profilePin_378 = core__GEN_388;
  wire  profilePin_379 = core__GEN_389;
  wire  profilePin_380 = core__GEN_390_0;
  wire  profilePin_381 = core__GEN_391;
  wire  profilePin_382 = core__GEN_392;
  wire  profilePin_383 = core__GEN_393_0;
  wire  profilePin_384 = core__GEN_394;
  wire  profilePin_385 = core__GEN_395;
  wire  profilePin_386 = core__GEN_396_0;
  wire [387:0] _GEN_1181 = {_GEN_1172,profilePin_378,profilePin_379,profilePin_380,profilePin_381,profilePin_382,profilePin_383,profilePin_384,profilePin_385,profilePin_386};
  wire  profilePin_387 = core__GEN_397;
  wire  profilePin_388 = core__GEN_398;
  wire  profilePin_389 = core__GEN_399_0;
  wire  profilePin_390 = core__GEN_400;
  wire  profilePin_391 = core__GEN_401;
  wire  profilePin_392 = core__GEN_402_0;
  wire  profilePin_393 = core__GEN_403;
  wire  profilePin_394 = core__GEN_404;
  wire  profilePin_395 = core__GEN_405_0;
  wire [396:0] _GEN_1190 = {_GEN_1181,profilePin_387,profilePin_388,profilePin_389,profilePin_390,profilePin_391,profilePin_392,profilePin_393,profilePin_394,profilePin_395};
  wire  profilePin_396 = core__GEN_406_0;
  wire  profilePin_397 = core__GEN_407;
  wire  profilePin_398 = core__GEN_408_0;
  wire  profilePin_399 = core__GEN_409_0;
  wire  profilePin_400 = core__GEN_410;
  wire  profilePin_401 = core__GEN_411;
  wire  profilePin_402 = core__GEN_412_0;
  wire  profilePin_403 = core__GEN_413;
  wire  profilePin_404 = core__GEN_414;
  wire [405:0] _GEN_1199 = {_GEN_1190,profilePin_396,profilePin_397,profilePin_398,profilePin_399,profilePin_400,profilePin_401,profilePin_402,profilePin_403,profilePin_404};
  wire  profilePin_405 = core__GEN_415_0;
  wire  profilePin_406 = core__GEN_416;
  wire  profilePin_407 = core__GEN_417;
  wire  profilePin_408 = core__GEN_418_0;
  wire  profilePin_409 = core__GEN_419;
  wire  profilePin_410 = core__GEN_420;
  wire  profilePin_411 = core__GEN_421;
  wire  profilePin_412 = core__GEN_422;
  wire  profilePin_413 = core__GEN_423;
  wire [414:0] _GEN_1208 = {_GEN_1199,profilePin_405,profilePin_406,profilePin_407,profilePin_408,profilePin_409,profilePin_410,profilePin_411,profilePin_412,profilePin_413};
  wire  profilePin_414 = core__GEN_424_0;
  wire  profilePin_415 = core__GEN_425;
  wire  profilePin_416 = core__GEN_0;
  wire  profilePin_417 = core__GEN_1_2;
  wire  profilePin_418 = core__GEN_3;
  wire  profilePin_419 = core__GEN_5_1;
  wire  profilePin_420 = core__GEN_6;
  wire  profilePin_421 = core__GEN_7;
  wire  profilePin_422 = core__GEN_11;
  wire [423:0] _GEN_1217 = {_GEN_1208,profilePin_414,profilePin_415,profilePin_416,profilePin_417,profilePin_418,profilePin_419,profilePin_420,profilePin_421,profilePin_422};
  wire  profilePin_423 = core__GEN_15_0;
  wire  profilePin_424 = core__GEN_146;
  wire  profilePin_425 = core__GEN_147_1;
  wire  profilePin_426 = core__GEN_149_0;
  wire  profilePin_427 = core__GEN_150;
  wire  profilePin_428 = core__GEN_151;
  wire  profilePin_429 = core__GEN_152_0;
  wire  profilePin_430 = core__GEN_234_0;
  wire  profilePin_431 = core__GEN_235_0;
  wire [432:0] _GEN_1226 = {_GEN_1217,profilePin_423,profilePin_424,profilePin_425,profilePin_426,profilePin_427,profilePin_428,profilePin_429,profilePin_430,profilePin_431};
  wire  profilePin_432 = core__GEN_236_0;
  wire  profilePin_433 = core__GEN_237;
  wire  profilePin_434 = core__GEN_238;
  wire  profilePin_435 = core__GEN_239_0;
  wire  profilePin_436 = core__GEN_240_0;
  wire  profilePin_437 = core__GEN_241_0;
  wire  profilePin_438 = core__GEN_242_0;
  wire  profilePin_439 = core__GEN_243;
  wire  profilePin_440 = core__GEN_244;
  wire [441:0] _GEN_1235 = {_GEN_1226,profilePin_432,profilePin_433,profilePin_434,profilePin_435,profilePin_436,profilePin_437,profilePin_438,profilePin_439,profilePin_440};
  wire  profilePin_441 = core__GEN_245_0;
  wire  profilePin_442 = core__GEN_246_0;
  wire  profilePin_443 = core__GEN_247_0;
  wire  profilePin_444 = core__GEN_248_0;
  wire  profilePin_445 = core__GEN_249_0;
  wire  profilePin_446 = core__GEN_250_0;
  wire  profilePin_447 = core__GEN_251_0;
  wire  profilePin_448 = core__GEN_252_0;
  wire  profilePin_449 = core__GEN_253;
  wire [450:0] _GEN_1244 = {_GEN_1235,profilePin_441,profilePin_442,profilePin_443,profilePin_444,profilePin_445,profilePin_446,profilePin_447,profilePin_448,profilePin_449};
  wire  profilePin_450 = core__GEN_254_0;
  wire  profilePin_451 = core__GEN_255;
  wire  profilePin_452 = core__GEN_256_0;
  wire  profilePin_453 = core__GEN_257_0;
  wire  profilePin_454 = core__GEN_258;
  wire  profilePin_455 = core__GEN_259_0;
  wire  profilePin_456 = core__GEN_260_0;
  wire  profilePin_457 = core__GEN_261;
  wire  profilePin_458 = core__GEN_262_0;
  wire [459:0] _GEN_1253 = {_GEN_1244,profilePin_450,profilePin_451,profilePin_452,profilePin_453,profilePin_454,profilePin_455,profilePin_456,profilePin_457,profilePin_458};
  wire  profilePin_459 = core__GEN_263_0;
  wire  profilePin_460 = core__GEN_264;
  wire  profilePin_461 = core__GEN_265_0;
  wire  profilePin_462 = core__GEN_266_0;
  wire  profilePin_463 = core__GEN_267_0;
  wire  profilePin_464 = core__GEN_268_0;
  wire  profilePin_465 = core__GEN_269_0;
  wire  profilePin_466 = core__GEN_270;
  wire  profilePin_467 = core__GEN_271_0;
  wire [468:0] _GEN_1262 = {_GEN_1253,profilePin_459,profilePin_460,profilePin_461,profilePin_462,profilePin_463,profilePin_464,profilePin_465,profilePin_466,profilePin_467};
  wire  profilePin_468 = core__GEN_272_0;
  wire  profilePin_469 = core__GEN_273;
  wire  profilePin_470 = core__GEN_274_0;
  wire  profilePin_471 = core__GEN_275_0;
  wire  profilePin_472 = core__GEN_276;
  wire  profilePin_473 = core__GEN_277_0;
  wire  profilePin_474 = core__GEN_278_0;
  wire  profilePin_475 = core__GEN_279;
  wire  profilePin_476 = core__GEN_280_0;
  wire [477:0] _GEN_1271 = {_GEN_1262,profilePin_468,profilePin_469,profilePin_470,profilePin_471,profilePin_472,profilePin_473,profilePin_474,profilePin_475,profilePin_476};
  wire  profilePin_477 = core__GEN_281_0;
  wire  profilePin_478 = core__GEN_282;
  wire  profilePin_479 = core__GEN_283_0;
  wire  profilePin_480 = core__GEN_284_0;
  wire  profilePin_481 = core__GEN_285;
  wire  profilePin_482 = core__GEN_286_0;
  wire  profilePin_483 = core__GEN_287_0;
  wire  profilePin_484 = core__GEN_288;
  wire  profilePin_485 = core__GEN_289_0;
  wire [486:0] _GEN_1280 = {_GEN_1271,profilePin_477,profilePin_478,profilePin_479,profilePin_480,profilePin_481,profilePin_482,profilePin_483,profilePin_484,profilePin_485};
  wire  profilePin_486 = core__GEN_290_0;
  wire  profilePin_487 = core__GEN_291;
  wire  profilePin_488 = core__GEN_292_0;
  wire  profilePin_489 = core__GEN_293_0;
  wire  profilePin_490 = core__GEN_294;
  wire  profilePin_491 = core__GEN_295_0;
  wire  profilePin_492 = core__GEN_296_0;
  wire  profilePin_493 = core__GEN_297;
  wire  profilePin_494 = core__GEN_298_0;
  wire [495:0] _GEN_1289 = {_GEN_1280,profilePin_486,profilePin_487,profilePin_488,profilePin_489,profilePin_490,profilePin_491,profilePin_492,profilePin_493,profilePin_494};
  wire  profilePin_495 = core__GEN_299_0;
  wire  profilePin_496 = core__GEN_300;
  wire  profilePin_497 = core__GEN_301_0;
  wire  profilePin_498 = core__GEN_302_0;
  wire  profilePin_499 = core__GEN_303;
  wire  profilePin_500 = core__GEN_304;
  wire  profilePin_501 = core__GEN_305_0;
  wire  profilePin_502 = core__GEN_306;
  wire  profilePin_503 = core__GEN_307;
  wire [504:0] _GEN_1298 = {_GEN_1289,profilePin_495,profilePin_496,profilePin_497,profilePin_498,profilePin_499,profilePin_500,profilePin_501,profilePin_502,profilePin_503};
  wire  profilePin_504 = core__GEN_308_0;
  wire  profilePin_505 = core__GEN_309;
  wire  profilePin_506 = core__GEN_310;
  wire  profilePin_507 = core__GEN_311_0;
  wire  profilePin_508 = core__GEN_312_0;
  wire  profilePin_509 = core__GEN_313;
  wire  profilePin_510 = core__GEN_314_0;
  wire  profilePin_511 = core__GEN_315_0;
  wire  profilePin_512 = core__GEN_316;
  wire [513:0] _GEN_1307 = {_GEN_1298,profilePin_504,profilePin_505,profilePin_506,profilePin_507,profilePin_508,profilePin_509,profilePin_510,profilePin_511,profilePin_512};
  wire  profilePin_513 = core__GEN_317_0;
  wire  profilePin_514 = core__GEN_318_0;
  wire  profilePin_515 = core__GEN_319;
  wire  profilePin_516 = core__GEN_320_0;
  wire  profilePin_517 = core__GEN_321_0;
  wire  profilePin_518 = core__GEN_322_0;
  wire  profilePin_519 = core__GEN_323_0;
  wire  profilePin_520 = core__GEN_324_0;
  wire  profilePin_521 = core__GEN_325;
  wire [522:0] _GEN_1316 = {_GEN_1307,profilePin_513,profilePin_514,profilePin_515,profilePin_516,profilePin_517,profilePin_518,profilePin_519,profilePin_520,profilePin_521};
  wire  profilePin_522 = core__GEN_326_0;
  wire  profilePin_523 = core__GEN_327_0;
  wire  profilePin_524 = core__GEN_328_0;
  wire  profilePin_525 = core__GEN_329_0;
  wire  profilePin_526 = core__GEN_330_0;
  wire  profilePin_527 = core__GEN_331;
  wire  profilePin_528 = core__GEN_332_0;
  wire  profilePin_529 = core__GEN_333_0;
  wire  profilePin_530 = core__GEN_334_0;
  wire [531:0] _GEN_1325 = {_GEN_1316,profilePin_522,profilePin_523,profilePin_524,profilePin_525,profilePin_526,profilePin_527,profilePin_528,profilePin_529,profilePin_530};
  wire  profilePin_531 = core__GEN_335_0;
  wire  profilePin_532 = core__GEN_336;
  wire  profilePin_533 = core__GEN_337;
  wire  profilePin_534 = core__GEN_338_0;
  wire  profilePin_535 = core__GEN_339_0;
  wire  profilePin_536 = core__GEN_340_0;
  wire  profilePin_537 = core__GEN_341_0;
  wire  profilePin_538 = core__GEN_342;
  wire  profilePin_539 = core__GEN_343_0;
  wire [540:0] _GEN_1334 = {_GEN_1325,profilePin_531,profilePin_532,profilePin_533,profilePin_534,profilePin_535,profilePin_536,profilePin_537,profilePin_538,profilePin_539};
  wire  profilePin_540 = core__GEN_344_0;
  wire  profilePin_541 = core__GEN_345_0;
  wire  profilePin_542 = core__GEN_346_0;
  wire  profilePin_543 = core__GEN_347_0;
  wire  profilePin_544 = core__GEN_348;
  wire  profilePin_545 = core__GEN_349_0;
  wire  profilePin_546 = core__GEN_350_0;
  wire  profilePin_547 = core__GEN_351_0;
  wire  profilePin_548 = core__GEN_352;
  wire [549:0] _GEN_1343 = {_GEN_1334,profilePin_540,profilePin_541,profilePin_542,profilePin_543,profilePin_544,profilePin_545,profilePin_546,profilePin_547,profilePin_548};
  wire  profilePin_549 = core__GEN_353_0;
  wire  profilePin_550 = core__GEN_354;
  wire  profilePin_551 = core__GEN_355_0;
  wire  profilePin_552 = core__GEN_356_0;
  wire  profilePin_553 = core__GEN_357;
  wire  profilePin_554 = core__GEN_358_0;
  wire  profilePin_555 = core__GEN_359_0;
  wire  profilePin_556 = core__GEN_360;
  wire  profilePin_557 = core__GEN_361_0;
  wire [558:0] _GEN_1352 = {_GEN_1343,profilePin_549,profilePin_550,profilePin_551,profilePin_552,profilePin_553,profilePin_554,profilePin_555,profilePin_556,profilePin_557};
  wire  profilePin_558 = core__GEN_362_0;
  wire  profilePin_559 = core__GEN_363;
  wire  profilePin_560 = core__GEN_364_0;
  wire  profilePin_561 = core__GEN_365_0;
  wire  profilePin_562 = core__GEN_366;
  wire  profilePin_563 = core__GEN_367_0;
  wire  profilePin_564 = core__GEN_368_0;
  wire  profilePin_565 = core__GEN_369;
  wire  profilePin_566 = core__GEN_370_0;
  wire [567:0] _GEN_1361 = {_GEN_1352,profilePin_558,profilePin_559,profilePin_560,profilePin_561,profilePin_562,profilePin_563,profilePin_564,profilePin_565,profilePin_566};
  wire  profilePin_567 = core__GEN_371_0;
  wire  profilePin_568 = core__GEN_372;
  wire  profilePin_569 = core__GEN_373_0;
  wire  profilePin_570 = core__GEN_374_0;
  wire  profilePin_571 = core__GEN_375;
  wire  profilePin_572 = core__GEN_376_0;
  wire  profilePin_573 = core__GEN_377_0;
  wire  profilePin_574 = core__GEN_378;
  wire  profilePin_575 = core__GEN_379_0;
  wire [576:0] _GEN_1370 = {_GEN_1361,profilePin_567,profilePin_568,profilePin_569,profilePin_570,profilePin_571,profilePin_572,profilePin_573,profilePin_574,profilePin_575};
  wire  profilePin_576 = core__GEN_380_0;
  wire  profilePin_577 = core__GEN_381;
  wire  profilePin_578 = core__GEN_382_0;
  wire  profilePin_579 = core__GEN_383_0;
  wire  profilePin_580 = core__GEN_384;
  wire  profilePin_581 = core__GEN_385_0;
  wire  profilePin_582 = core__GEN_386_0;
  wire  profilePin_583 = core__GEN_387;
  wire  profilePin_584 = core__GEN_388_0;
  wire [585:0] _GEN_1379 = {_GEN_1370,profilePin_576,profilePin_577,profilePin_578,profilePin_579,profilePin_580,profilePin_581,profilePin_582,profilePin_583,profilePin_584};
  wire  profilePin_585 = core__GEN_389_0;
  wire  profilePin_586 = core__GEN_390;
  wire  profilePin_587 = core__GEN_391_0;
  wire  profilePin_588 = core__GEN_392_0;
  wire  profilePin_589 = core__GEN_393;
  wire  profilePin_590 = core__GEN_394_0;
  wire  profilePin_591 = core__GEN_395_0;
  wire  profilePin_592 = core__GEN_396;
  wire  profilePin_593 = core__GEN_397_0;
  wire [594:0] _GEN_1388 = {_GEN_1379,profilePin_585,profilePin_586,profilePin_587,profilePin_588,profilePin_589,profilePin_590,profilePin_591,profilePin_592,profilePin_593};
  wire  profilePin_594 = core__GEN_398_0;
  wire  profilePin_595 = core__GEN_399;
  wire  profilePin_596 = core__GEN_400_0;
  wire  profilePin_597 = core__GEN_401_0;
  wire  profilePin_598 = core__GEN_402;
  wire  profilePin_599 = core__GEN_403_0;
  wire  profilePin_600 = core__GEN_404_0;
  wire  profilePin_601 = core__GEN_405;
  wire  profilePin_602 = core__GEN_406;
  wire [603:0] _GEN_1397 = {_GEN_1388,profilePin_594,profilePin_595,profilePin_596,profilePin_597,profilePin_598,profilePin_599,profilePin_600,profilePin_601,profilePin_602};
  wire  profilePin_603 = core__GEN_407_0;
  wire  profilePin_604 = core__GEN_408;
  wire  profilePin_605 = core__GEN_409;
  wire  profilePin_606 = core__GEN_410_0;
  wire  profilePin_607 = core__GEN_411_0;
  wire  profilePin_608 = core__GEN_412;
  wire  profilePin_609 = core__GEN_413_0;
  wire  profilePin_610 = core__GEN_414_0;
  wire  profilePin_611 = core__GEN_415;
  wire [612:0] _GEN_1406 = {_GEN_1397,profilePin_603,profilePin_604,profilePin_605,profilePin_606,profilePin_607,profilePin_608,profilePin_609,profilePin_610,profilePin_611};
  wire  profilePin_612 = core__GEN_416_0;
  wire  profilePin_613 = core__GEN_417_0;
  wire  profilePin_614 = core__GEN_418;
  wire  profilePin_615 = core__GEN_419_0;
  wire  profilePin_616 = core__GEN_420_0;
  wire  profilePin_617 = core__GEN_421_0;
  wire  profilePin_618 = core__GEN_422_0;
  wire  profilePin_619 = core__GEN_423_0;
  wire  profilePin_620 = core__GEN_424;
  wire [621:0] _GEN_1415 = {_GEN_1406,profilePin_612,profilePin_613,profilePin_614,profilePin_615,profilePin_616,profilePin_617,profilePin_618,profilePin_619,profilePin_620};
  wire  profilePin_621 = core__GEN_425_0;
  wire  profilePin_622 = core__GEN_426;
  wire  profilePin_623 = core__GEN_427;
  wire  profilePin_624 = core__GEN_428;
  wire  profilePin_625 = core__GEN_429;
  wire  profilePin_626 = core__GEN_430;
  wire  profilePin_627 = core__GEN_431;
  wire  profilePin_628 = core__GEN_432;
  wire  profilePin_629 = core__GEN_433;
  wire [630:0] _GEN_1424 = {_GEN_1415,profilePin_621,profilePin_622,profilePin_623,profilePin_624,profilePin_625,profilePin_626,profilePin_627,profilePin_628,profilePin_629};
  wire  profilePin_630 = core__GEN_434;
  wire  profilePin_631 = core__GEN_435;
  wire  profilePin_632 = core__GEN_436;
  wire  profilePin_633 = core__GEN_437;
  wire  profilePin_634 = core__GEN_438;
  wire  profilePin_635 = core__GEN_439;
  wire  profilePin_636 = core__GEN_440;
  wire  profilePin_637 = core__GEN_441;
  wire  profilePin_638 = core__GEN_442;
  wire [639:0] _GEN_1433 = {_GEN_1424,profilePin_630,profilePin_631,profilePin_632,profilePin_633,profilePin_634,profilePin_635,profilePin_636,profilePin_637,profilePin_638};
  wire  profilePin_639 = core__GEN_443;
  wire  profilePin_640 = core__GEN_444;
  wire  profilePin_641 = core__GEN_445;
  wire  profilePin_642 = core__GEN_446;
  wire  profilePin_643 = core__GEN_447;
  wire  profilePin_644 = core__GEN_448;
  wire  profilePin_645 = core__GEN_449;
  wire  profilePin_646 = core__GEN_450;
  wire  profilePin_647 = core__GEN_451;
  wire [648:0] _GEN_1442 = {_GEN_1433,profilePin_639,profilePin_640,profilePin_641,profilePin_642,profilePin_643,profilePin_644,profilePin_645,profilePin_646,profilePin_647};
  wire  profilePin_648 = core__GEN_452;
  wire  profilePin_649 = core__GEN_453;
  wire  profilePin_650 = core__GEN_454;
  wire  profilePin_651 = core__GEN_455;
  wire  profilePin_652 = core__GEN_456;
  wire  profilePin_653 = core__GEN_457;
  wire  profilePin_654 = core__GEN_458;
  wire  profilePin_655 = core__GEN_459;
  wire  profilePin_656 = core__GEN_460;
  wire [657:0] _GEN_1451 = {_GEN_1442,profilePin_648,profilePin_649,profilePin_650,profilePin_651,profilePin_652,profilePin_653,profilePin_654,profilePin_655,profilePin_656};
  wire  profilePin_657 = core__GEN_461;
  wire  profilePin_658 = core__GEN_462;
  wire  profilePin_660 = core__GEN_1_1;
  wire  profilePin_661 = core__GEN_16;
  wire  profilePin_662 = core__GEN_17_0;
  wire  profilePin_663 = core__GEN_21;
  wire  profilePin_664 = core__GEN_33;
  wire  profilePin_665 = core__GEN_40_0;
  wire  profilePin_666 = core__GEN_41_0;
  wire [666:0] _GEN_1460 = {_GEN_1451,profilePin_657,profilePin_658,profilePin_660,profilePin_661,profilePin_662,profilePin_663,profilePin_664,profilePin_665,profilePin_666};
  wire  profilePin_667 = core__GEN_42;
  wire  profilePin_668 = core__GEN_43_0;
  wire  profilePin_669 = core__GEN_44_0;
  wire  profilePin_670 = core__GEN_45;
  wire  profilePin_671 = core__GEN_46_0;
  wire  profilePin_672 = core__GEN_47_0;
  wire  profilePin_673 = core__GEN_53_0;
  wire  profilePin_674 = core__GEN_54_0;
  wire  profilePin_675 = core__GEN_55_0;
  wire [675:0] _GEN_1469 = {_GEN_1460,profilePin_667,profilePin_668,profilePin_669,profilePin_670,profilePin_671,profilePin_672,profilePin_673,profilePin_674,profilePin_675};
  wire  profilePin_676 = core__GEN_56;
  wire  profilePin_677 = core__GEN_64_0;
  wire  profilePin_678 = core__GEN_68_0;
  wire  profilePin_679 = core__GEN_69;
  wire  profilePin_680 = core__GEN_70_0;
  wire  profilePin_681 = core__GEN_71_0;
  wire  profilePin_682 = core__GEN_72;
  wire  profilePin_683 = core__GEN_73_0;
  wire  profilePin_684 = core__GEN_74_0;
  wire [684:0] _GEN_1478 = {_GEN_1469,profilePin_676,profilePin_677,profilePin_678,profilePin_679,profilePin_680,profilePin_681,profilePin_682,profilePin_683,profilePin_684};
  wire  profilePin_685 = core__GEN_75;
  wire  profilePin_686 = core__GEN_78_0;
  wire  profilePin_687 = core__GEN_79;
  wire  profilePin_688 = core__GEN_80;
  wire  profilePin_689 = core__GEN_82_0;
  wire  profilePin_690 = core__GEN_83;
  wire  profilePin_691 = core__GEN_85;
  wire  profilePin_692 = core__GEN_86_0;
  wire  profilePin_693 = core__GEN_87;
  wire [693:0] _GEN_1487 = {_GEN_1478,profilePin_685,profilePin_686,profilePin_687,profilePin_688,profilePin_689,profilePin_690,profilePin_691,profilePin_692,profilePin_693};
  wire  profilePin_694 = core__GEN_88;
  wire  profilePin_695 = core__GEN_89;
  wire  profilePin_696 = core__GEN_90;
  wire  profilePin_697 = core__GEN_91;
  wire  profilePin_698 = core__GEN_92_0;
  wire  profilePin_699 = core__GEN_93;
  wire  profilePin_700 = core__GEN_94_0;
  wire  profilePin_701 = core__GEN_95;
  wire  profilePin_702 = core__GEN_96_0;
  wire [702:0] _GEN_1496 = {_GEN_1487,profilePin_694,profilePin_695,profilePin_696,profilePin_697,profilePin_698,profilePin_699,profilePin_700,profilePin_701,profilePin_702};
  wire  profilePin_703 = core__GEN_97_0;
  wire  profilePin_704 = core__GEN_98;
  wire  profilePin_705 = core__GEN_99_0;
  wire  profilePin_706 = core__GEN_100_0;
  wire  profilePin_707 = core__GEN_101;
  wire  profilePin_708 = core__GEN_102_0;
  wire  profilePin_709 = core__GEN_103;
  wire  profilePin_710 = core__GEN_104;
  wire  profilePin_711 = core__GEN_105_0;
  wire [711:0] _GEN_1505 = {_GEN_1496,profilePin_703,profilePin_704,profilePin_705,profilePin_706,profilePin_707,profilePin_708,profilePin_709,profilePin_710,profilePin_711};
  wire  profilePin_712 = core__GEN_106_0;
  wire  profilePin_713 = core__GEN_107;
  wire  profilePin_714 = core__GEN_108_0;
  wire  profilePin_715 = core__GEN_109_0;
  wire  profilePin_716 = core__GEN_110_0;
  wire  profilePin_717 = core__GEN_111_0;
  wire  profilePin_718 = core__GEN_112;
  wire  profilePin_719 = core__GEN_113;
  wire  profilePin_720 = core__GEN_114_0;
  wire [720:0] _GEN_1514 = {_GEN_1505,profilePin_712,profilePin_713,profilePin_714,profilePin_715,profilePin_716,profilePin_717,profilePin_718,profilePin_719,profilePin_720};
  wire  profilePin_721 = core__GEN_115;
  wire  profilePin_722 = core__GEN_116_0;
  wire  profilePin_723 = core__GEN_117_0;
  wire  profilePin_724 = core__GEN_118;
  wire  profilePin_725 = core__GEN_119;
  wire  profilePin_726 = core__GEN_120_0;
  wire  profilePin_727 = core__GEN_121;
  wire  profilePin_728 = core__GEN_122;
  wire  profilePin_729 = core__GEN_123_0;
  wire [729:0] _GEN_1523 = {_GEN_1514,profilePin_721,profilePin_722,profilePin_723,profilePin_724,profilePin_725,profilePin_726,profilePin_727,profilePin_728,profilePin_729};
  wire  profilePin_730 = core__GEN_124;
  wire  profilePin_731 = core__GEN_125;
  wire  profilePin_732 = core__GEN_126_0;
  wire  profilePin_733 = core__GEN_127;
  wire  profilePin_734 = core__GEN_128_0;
  wire  profilePin_735 = core__GEN_129_0;
  wire  profilePin_736 = core__GEN_130;
  wire  profilePin_737 = core__GEN_131_0;
  wire  profilePin_738 = core__GEN_132_0;
  wire [738:0] _GEN_1532 = {_GEN_1523,profilePin_730,profilePin_731,profilePin_732,profilePin_733,profilePin_734,profilePin_735,profilePin_736,profilePin_737,profilePin_738};
  wire  profilePin_739 = core__GEN_133;
  wire  profilePin_740 = core__GEN_134_0;
  wire  profilePin_741 = core__GEN_135_0;
  wire  profilePin_742 = core__GEN_136;
  wire  profilePin_743 = core__GEN_137_0;
  wire  profilePin_744 = core__GEN_138;
  wire  profilePin_745 = core__GEN_139;
  wire  profilePin_746 = core__GEN_140;
  wire  profilePin_747 = core__GEN_141_0;
  wire [747:0] _GEN_1541 = {_GEN_1532,profilePin_739,profilePin_740,profilePin_741,profilePin_742,profilePin_743,profilePin_744,profilePin_745,profilePin_746,profilePin_747};
  wire  profilePin_748 = core__GEN_142;
  wire  profilePin_749 = core__GEN_143_0;
  wire  profilePin_750 = core__GEN_144;
  wire  profilePin_751 = core__GEN_145;
  wire  profilePin_752 = core__GEN_146_1;
  wire  profilePin_753 = core__GEN_147_0;
  wire  profilePin_754 = core__GEN_148;
  wire  profilePin_755 = core__GEN_149_1;
  wire  profilePin_756 = core__GEN_150_0;
  wire [756:0] _GEN_1550 = {_GEN_1541,profilePin_748,profilePin_749,profilePin_750,profilePin_751,profilePin_752,profilePin_753,profilePin_754,profilePin_755,profilePin_756};
  wire  profilePin_757 = core__GEN_151_0;
  wire  profilePin_758 = core__GEN_152_1;
  wire  profilePin_759 = core__GEN_153_0;
  wire  profilePin_760 = core__GEN_154;
  wire  profilePin_761 = core__GEN_155_0;
  wire  profilePin_762 = core__GEN_156;
  wire  profilePin_763 = core__GEN_157;
  wire  profilePin_764 = core__GEN_158_0;
  wire  profilePin_765 = core__GEN_159;
  wire [765:0] _GEN_1559 = {_GEN_1550,profilePin_757,profilePin_758,profilePin_759,profilePin_760,profilePin_761,profilePin_762,profilePin_763,profilePin_764,profilePin_765};
  wire  profilePin_766 = core__GEN_160;
  wire  profilePin_767 = core__GEN_161_0;
  wire  profilePin_768 = core__GEN_162;
  wire  profilePin_769 = core__GEN_163;
  wire  profilePin_770 = core__GEN_164_0;
  wire  profilePin_771 = core__GEN_165;
  wire  profilePin_772 = core__GEN_166;
  wire  profilePin_773 = core__GEN_167_0;
  wire  profilePin_774 = core__GEN_168_0;
  wire [774:0] _GEN_1568 = {_GEN_1559,profilePin_766,profilePin_767,profilePin_768,profilePin_769,profilePin_770,profilePin_771,profilePin_772,profilePin_773,profilePin_774};
  wire  profilePin_775 = core__GEN_169;
  wire  profilePin_776 = core__GEN_170_0;
  wire  profilePin_777 = core__GEN_171;
  wire  profilePin_778 = core__GEN_172;
  wire  profilePin_779 = core__GEN_173_0;
  wire  profilePin_780 = core__GEN_174;
  wire  profilePin_781 = core__GEN_175;
  wire  profilePin_782 = core__GEN_176_0;
  wire  profilePin_783 = core__GEN_177;
  wire [783:0] _GEN_1577 = {_GEN_1568,profilePin_775,profilePin_776,profilePin_777,profilePin_778,profilePin_779,profilePin_780,profilePin_781,profilePin_782,profilePin_783};
  wire  profilePin_784 = core__GEN_178;
  wire  profilePin_785 = core__GEN_179_0;
  wire  profilePin_786 = memory__GEN_0_1;
  wire  profilePin_787 = memory__GEN_1_1;
  wire  profilePin_788 = memory__GEN_2_0;
  wire  profilePin_789 = memory__GEN_3_1;
  wire  profilePin_790 = memory__GEN_4_0;
  wire [790:0] _GEN_1584 = {_GEN_1577,profilePin_784,profilePin_785,profilePin_786,profilePin_787,profilePin_788,profilePin_789,profilePin_790};
  wire  profilePin_791 = memory__GEN_5_0;
  Core core ( // @[top.scala 21:26]
    .metaReset(core_metaReset),
    .clock(core_clock),
    .reset(core_reset),
    .io_imem_req_bits_addr(core_io_imem_req_bits_addr),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_imem_resp_bits_data(core_io_imem_resp_bits_data),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_data(core_io_dmem_req_bits_data),
    .io_dmem_req_bits_fcn(core_io_dmem_req_bits_fcn),
    .io_dmem_req_bits_typ(core_io_dmem_req_bits_typ),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
    ._GEN_451(core__GEN_451),
    ._GEN_331(core__GEN_331),
    ._GEN_337(core__GEN_337),
    ._GEN_113(core__GEN_113),
    ._GEN_111(core__GEN_111),
    ._GEN_415(core__GEN_415),
    ._GEN_436(core__GEN_436),
    ._GEN_140(core__GEN_140),
    ._GEN_71(core__GEN_71),
    ._GEN_324(core__GEN_324),
    ._GEN_219(core__GEN_219),
    ._GEN_168(core__GEN_168),
    ._GEN_98(core__GEN_98),
    ._GEN_1(core__GEN_1),
    ._GEN_352(core__GEN_352),
    ._GEN_423(core__GEN_423),
    ._GEN_44(core__GEN_44),
    ._GEN_125(core__GEN_125),
    ._GEN_267(core__GEN_267),
    ._GEN_126(core__GEN_126),
    ._GEN_430(core__GEN_430),
    ._GEN_153(core__GEN_153),
    ._GEN_225(core__GEN_225),
    ._GEN_119(core__GEN_119),
    ._GEN_88(core__GEN_88),
    ._GEN_59(core__GEN_59),
    ._GEN_252(core__GEN_252),
    ._GEN_151(core__GEN_151),
    ._GEN_147(core__GEN_147),
    ._GEN_310(core__GEN_310),
    ._GEN_351(core__GEN_351),
    ._GEN_210(core__GEN_210),
    ._GEN_246(core__GEN_246),
    ._GEN_104(core__GEN_104),
    ._GEN_409(core__GEN_409),
    ._GEN_65(core__GEN_65),
    ._GEN_253(core__GEN_253),
    ._GEN_132(core__GEN_132),
    ._GEN_318(core__GEN_318),
    ._GEN_316(core__GEN_316),
    ._GEN_92(core__GEN_92),
    ._GEN_345(core__GEN_345),
    ._GEN_231(core__GEN_231),
    ._GEN_417(core__GEN_417),
    ._GEN_244(core__GEN_244),
    ._GEN_50(core__GEN_50),
    ._GEN_238(core__GEN_238),
    ._GEN_330(core__GEN_330),
    ._GEN_86(core__GEN_86),
    ._GEN_339(core__GEN_339),
    ._GEN_101(core__GEN_101),
    ._GEN_325(core__GEN_325),
    ._GEN_240(core__GEN_240),
    ._GEN_234(core__GEN_234),
    ._GEN_120(core__GEN_120),
    ._GEN_169(core__GEN_169),
    ._GEN_129(core__GEN_129),
    ._GEN_433(core__GEN_433),
    ._GEN_333(core__GEN_333),
    ._GEN_302(core__GEN_302),
    ._GEN_313(core__GEN_313),
    ._GEN_228(core__GEN_228),
    ._GEN_197(core__GEN_197),
    ._GEN_91(core__GEN_91),
    ._GEN_411(core__GEN_411),
    ._GEN_11(core__GEN_11),
    ._GEN_401(core__GEN_401),
    ._GEN_47(core__GEN_47),
    ._GEN_296(core__GEN_296),
    ._GEN_304(core__GEN_304),
    ._GEN_294(core__GEN_294),
    ._GEN_74(core__GEN_74),
    ._GEN_213(core__GEN_213),
    ._GEN_303(core__GEN_303),
    ._GEN_107(core__GEN_107),
    ._GEN_32(core__GEN_32),
    ._GEN_0(core__GEN_0),
    ._GEN_402(core__GEN_402),
    ._GEN_412(core__GEN_412),
    ._GEN_68(core__GEN_68),
    ._GEN_135(core__GEN_135),
    ._GEN_424(core__GEN_424),
    ._GEN_175(core__GEN_175),
    ._GEN_319(core__GEN_319),
    ._GEN_288(core__GEN_288),
    ._GEN_56(core__GEN_56),
    ._GEN_26(core__GEN_26),
    ._GEN_418(core__GEN_418),
    ._GEN_122(core__GEN_122),
    ._GEN_387(core__GEN_387),
    ._GEN_53(core__GEN_53),
    ._GEN_141(core__GEN_141),
    ._GEN_327(core__GEN_327),
    ._GEN_72(core__GEN_72),
    ._GEN_395(core__GEN_395),
    ._GEN_249(core__GEN_249),
    ._GEN_114(core__GEN_114),
    ._GEN_312(core__GEN_312),
    ._GEN_203(core__GEN_203),
    ._GEN_75(core__GEN_75),
    ._GEN_85(core__GEN_85),
    ._GEN_20(core__GEN_20),
    ._GEN_178(core__GEN_178),
    ._GEN_15(core__GEN_15),
    ._GEN_157(core__GEN_157),
    ._GEN_462(core__GEN_462),
    ._GEN_69(core__GEN_69),
    ._GEN_216(core__GEN_216),
    ._GEN_206(core__GEN_206),
    ._GEN_375(core__GEN_375),
    ._GEN_151_0(core__GEN_151_0),
    ._GEN_420(core__GEN_420),
    ._GEN_123(core__GEN_123),
    ._GEN_315(core__GEN_315),
    ._GEN_284(core__GEN_284),
    ._GEN_179(core__GEN_179),
    ._GEN_33(core__GEN_33),
    ._GEN_222(core__GEN_222),
    ._GEN_377(core__GEN_377),
    ._GEN_191(core__GEN_191),
    ._GEN_290(core__GEN_290),
    ._GEN_404(core__GEN_404),
    ._GEN_390(core__GEN_390),
    ._GEN_56_0(core__GEN_56_0),
    ._GEN_305(core__GEN_305),
    ._GEN_299(core__GEN_299),
    ._GEN_185(core__GEN_185),
    ._GEN_307(core__GEN_307),
    ._GEN_297(core__GEN_297),
    ._GEN_398(core__GEN_398),
    ._GEN_406(core__GEN_406),
    ._GEN_41(core__GEN_41),
    ._GEN_321(core__GEN_321),
    ._GEN_270(core__GEN_270),
    ._GEN_95(core__GEN_95),
    ._GEN_45(core__GEN_45),
    ._GEN_414(core__GEN_414),
    ._GEN_383(core__GEN_383),
    ._GEN_369(core__GEN_369),
    ._GEN_35(core__GEN_35),
    ._GEN_29(core__GEN_29),
    ._GEN_278(core__GEN_278),
    ._GEN_117(core__GEN_117),
    ._GEN_396(core__GEN_396),
    ._GEN_172(core__GEN_172),
    ._GEN_276(core__GEN_276),
    ._GEN_291(core__GEN_291),
    ._GEN_365(core__GEN_365),
    ._GEN_359(core__GEN_359),
    ._GEN_258(core__GEN_258),
    ._GEN_372(core__GEN_372),
    ._GEN_38(core__GEN_38),
    ._GEN_252_0(core__GEN_252_0),
    ._GEN_167(core__GEN_167),
    ._GEN_166(core__GEN_166),
    ._GEN_285(core__GEN_285),
    ._GEN_42(core__GEN_42),
    ._GEN_350(core__GEN_350),
    ._GEN_106(core__GEN_106),
    ._GEN_384(core__GEN_384),
    ._GEN_18(core__GEN_18),
    ._GEN_378(core__GEN_378),
    ._GEN_393(core__GEN_393),
    ._GEN_273(core__GEN_273),
    ._GEN_293(core__GEN_293),
    ._GEN_456(core__GEN_456),
    ._GEN_371(core__GEN_371),
    ._GEN_80(core__GEN_80),
    ._GEN_351_0(core__GEN_351_0),
    ._GEN_251(core__GEN_251),
    ._GEN_209(core__GEN_209),
    ._GEN_139(core__GEN_139),
    ._GEN_145(core__GEN_145),
    ._GEN_450(core__GEN_450),
    ._GEN_308(core__GEN_308),
    ._GEN_173(core__GEN_173),
    ._GEN_53_0(core__GEN_53_0),
    ._GEN_357(core__GEN_357),
    ._GEN_200(core__GEN_200),
    ._GEN_386(core__GEN_386),
    ._GEN_272(core__GEN_272),
    ._GEN_160(core__GEN_160),
    ._GEN_91_0(core__GEN_91_0),
    ._GEN_279(core__GEN_279),
    ._GEN_194(core__GEN_194),
    ._GEN_188(core__GEN_188),
    ._GEN_133(core__GEN_133),
    ._GEN_392(core__GEN_392),
    ._GEN_23(core__GEN_23),
    ._GEN_407(core__GEN_407),
    ._GEN_287(core__GEN_287),
    ._GEN_266(core__GEN_266),
    ._GEN_399(core__GEN_399),
    ._GEN_264(core__GEN_264),
    ._GEN_300(core__GEN_300),
    ._GEN_374(core__GEN_374),
    ._GEN_233(core__GEN_233),
    ._GEN_127(core__GEN_127),
    ._GEN_269(core__GEN_269),
    ._GEN_432(core__GEN_432),
    ._GEN_381(core__GEN_381),
    ._GEN_260(core__GEN_260),
    ._GEN_161(core__GEN_161),
    ._GEN_155(core__GEN_155),
    ._GEN_339_0(core__GEN_339_0),
    ._GEN_368(core__GEN_368),
    ._GEN_254(core__GEN_254),
    ._GEN_281(core__GEN_281),
    ._GEN_73(core__GEN_73),
    ._GEN_261(core__GEN_261),
    ._GEN_353(core__GEN_353),
    ._GEN_332(core__GEN_332),
    ._GEN_88_0(core__GEN_88_0),
    ._GEN_176(core__GEN_176),
    ._GEN_16(core__GEN_16),
    ._GEN_380(core__GEN_380),
    ._GEN_360(core__GEN_360),
    ._GEN_389(core__GEN_389),
    ._GEN_163(core__GEN_163),
    ._GEN_246_0(core__GEN_246_0),
    ._GEN_438(core__GEN_438),
    ._GEN_94(core__GEN_94),
    ._GEN_282(core__GEN_282),
    ._GEN_347(core__GEN_347),
    ._GEN_109(core__GEN_109),
    ._GEN_182(core__GEN_182),
    ._GEN_345_0(core__GEN_345_0),
    ._GEN_121(core__GEN_121),
    ._GEN_240_0(core__GEN_240_0),
    ._GEN_9(core__GEN_9),
    ._GEN_148(core__GEN_148),
    ._GEN_154(core__GEN_154),
    ._GEN_444(core__GEN_444),
    ._GEN_149(core__GEN_149),
    ._GEN_267_0(core__GEN_267_0),
    ._GEN_459(core__GEN_459),
    ._GEN_453(core__GEN_453),
    ._GEN_248(core__GEN_248),
    ._GEN_366(core__GEN_366),
    ._GEN_7(core__GEN_7),
    ._GEN_142(core__GEN_142),
    ._GEN_275(core__GEN_275),
    ._GEN_140_0(core__GEN_140_0),
    ._GEN_324_0(core__GEN_324_0),
    ._GEN_100(core__GEN_100),
    ._GEN_333_0(core__GEN_333_0),
    ._GEN_362(core__GEN_362),
    ._GEN_413(core__GEN_413),
    ._GEN_342(core__GEN_342),
    ._GEN_405(core__GEN_405),
    ._GEN_420_0(core__GEN_420_0),
    ._GEN_306(core__GEN_306),
    ._GEN_76(core__GEN_76),
    ._GEN_164(core__GEN_164),
    ._GEN_109_0(core__GEN_109_0),
    ._GEN_103(core__GEN_103),
    ._GEN_3(core__GEN_3),
    ._GEN_242(core__GEN_242),
    ._GEN_136(core__GEN_136),
    ._GEN_426(core__GEN_426),
    ._GEN_137(core__GEN_137),
    ._GEN_441(core__GEN_441),
    ._GEN_341(core__GEN_341),
    ._GEN_94_0(core__GEN_94_0),
    ._GEN_348(core__GEN_348),
    ._GEN_263(core__GEN_263),
    ._GEN_257(core__GEN_257),
    ._GEN_122_0(core__GEN_122_0),
    ._GEN_143(core__GEN_143),
    ._GEN_255(core__GEN_255),
    ._GEN_82(core__GEN_82),
    ._GEN_170(core__GEN_170),
    ._GEN_356(core__GEN_356),
    ._GEN_221(core__GEN_221),
    ._GEN_215(core__GEN_215),
    ._GEN_115(core__GEN_115),
    ._GEN_146(core__GEN_146),
    ._GEN_363(core__GEN_363),
    ._GEN_320(core__GEN_320),
    ._GEN_314(core__GEN_314),
    ._GEN_329(core__GEN_329),
    ._GEN_321_0(core__GEN_321_0),
    ._GEN_327_0(core__GEN_327_0),
    ._GEN_103_0(core__GEN_103_0),
    ._GEN_97(core__GEN_97),
    ._GEN_236(core__GEN_236),
    ._GEN_354(core__GEN_354),
    ._GEN_234_0(core__GEN_234_0),
    ._GEN_130(core__GEN_130),
    ._GEN_61(core__GEN_61),
    ._GEN_55(core__GEN_55),
    ._GEN_249_0(core__GEN_249_0),
    ._GEN_335(core__GEN_335),
    ._GEN_243(core__GEN_243),
    ._GEN_447(core__GEN_447),
    ._GEN_158(core__GEN_158),
    ._GEN_330_0(core__GEN_330_0),
    ._GEN_422(core__GEN_422),
    ._GEN_245(core__GEN_245),
    ._GEN_37(core__GEN_37),
    ._GEN_125_0(core__GEN_125_0),
    ._GEN_429(core__GEN_429),
    ._GEN_70(core__GEN_70),
    ._GEN_64(core__GEN_64),
    ._GEN_344(core__GEN_344),
    ._GEN_338(core__GEN_338),
    ._GEN_293_0(core__GEN_293_0),
    ._GEN_87(core__GEN_87),
    ._GEN_416(core__GEN_416),
    ._GEN_406_0(core__GEN_406_0),
    ._GEN_58(core__GEN_58),
    ._GEN_414_0(core__GEN_414_0),
    ._GEN_309(core__GEN_309),
    ._GEN_85_0(core__GEN_85_0),
    ._GEN_299_0(core__GEN_299_0),
    ._GEN_336(core__GEN_336),
    ._GEN_408(core__GEN_408),
    ._GEN_112(core__GEN_112),
    ._GEN_43(core__GEN_43),
    ._GEN_150(core__GEN_150),
    ._GEN_131(core__GEN_131),
    ._GEN_435(core__GEN_435),
    ._GEN_230(core__GEN_230),
    ._GEN_97_0(core__GEN_97_0),
    ._GEN_124(core__GEN_124),
    ._GEN_239(core__GEN_239),
    ._GEN_118(core__GEN_118),
    ._GEN_392_0(core__GEN_392_0),
    ._GEN_398_0(core__GEN_398_0),
    ._GEN_423_0(core__GEN_423_0),
    ._GEN_237(core__GEN_237),
    ._GEN_152(core__GEN_152),
    ._GEN_307_0(core__GEN_307_0),
    ._GEN_146_0(core__GEN_146_0),
    ._GEN_315_0(core__GEN_315_0),
    ._GEN_79(core__GEN_79),
    ._GEN_224(core__GEN_224),
    ._GEN_110(core__GEN_110),
    ._GEN_119_0(core__GEN_119_0),
    ._GEN_323(core__GEN_323),
    ._GEN_317(core__GEN_317),
    ._GEN_79_0(core__GEN_79_0),
    ._GEN_218(core__GEN_218),
    ._GEN_208(core__GEN_208),
    ._GEN_1_1(core__GEN_1_1),
    ._GEN_196(core__GEN_196),
    ._GEN_90(core__GEN_90),
    ._GEN_31(core__GEN_31),
    ._GEN_400(core__GEN_400),
    ._GEN_113_0(core__GEN_113_0),
    ._GEN_162(core__GEN_162),
    ._GEN_212(core__GEN_212),
    ._GEN_302_0(core__GEN_302_0),
    ._GEN_181(core__GEN_181),
    ._GEN_106_0(core__GEN_106_0),
    ._GEN_227(core__GEN_227),
    ._GEN_71_0(core__GEN_71_0),
    ._GEN_380_0(core__GEN_380_0),
    ._GEN_425(core__GEN_425),
    ._GEN_280(core__GEN_280),
    ._GEN_46(core__GEN_46),
    ._GEN_174(core__GEN_174),
    ._GEN_134(core__GEN_134),
    ._GEN_289(core__GEN_289),
    ._GEN_318_0(core__GEN_318_0),
    ._GEN_287_0(core__GEN_287_0),
    ._GEN_202(core__GEN_202),
    ._GEN_419(core__GEN_419),
    ._GEN_388(core__GEN_388),
    ._GEN_410(core__GEN_410),
    ._GEN_386_0(core__GEN_386_0),
    ._GEN_52(core__GEN_52),
    ._GEN_311(core__GEN_311),
    ._GEN_301(core__GEN_301),
    ._GEN_295(core__GEN_295),
    ._GEN_67(core__GEN_67),
    ._GEN_281_0(core__GEN_281_0),
    ._GEN_312_0(core__GEN_312_0),
    ._GEN_25(core__GEN_25),
    ._GEN_409_0(core__GEN_409_0),
    ._GEN_417_0(core__GEN_417_0),
    ._GEN_411_0(core__GEN_411_0),
    ._GEN_326(core__GEN_326),
    ._GEN_55_0(core__GEN_55_0),
    ._GEN_100_0(core__GEN_100_0),
    ._GEN_394(core__GEN_394),
    ._GEN_168_0(core__GEN_168_0),
    ._GEN_128(core__GEN_128),
    ._GEN_401_0(core__GEN_401_0),
    ._GEN_44_0(core__GEN_44_0),
    ._GEN_376(core__GEN_376),
    ._GEN_74_0(core__GEN_74_0),
    ._GEN_374_0(core__GEN_374_0),
    ._GEN_40(core__GEN_40),
    ._GEN_368_0(core__GEN_368_0),
    ._GEN_34(core__GEN_34),
    ._GEN_383_0(core__GEN_383_0),
    ._GEN_49(core__GEN_49),
    ._GEN_263_0(core__GEN_263_0),
    ._GEN_177(core__GEN_177),
    ._GEN_171(core__GEN_171),
    ._GEN_446(core__GEN_446),
    ._GEN_102(core__GEN_102),
    ._GEN_290_0(core__GEN_290_0),
    ._GEN_190(core__GEN_190),
    ._GEN_83(core__GEN_83),
    ._GEN_205(core__GEN_205),
    ._GEN_135_0(core__GEN_135_0),
    ._GEN_389_0(core__GEN_389_0),
    ._GEN_93(core__GEN_93),
    ._GEN_254_0(core__GEN_254_0),
    ._GEN_298(core__GEN_298),
    ._GEN_163_0(core__GEN_163_0),
    ._GEN_21(core__GEN_21),
    ._GEN_461(core__GEN_461),
    ._GEN_362_0(core__GEN_362_0),
    ._GEN_14(core__GEN_14),
    ._GEN_116(core__GEN_116),
    ._GEN_156(core__GEN_156),
    ._GEN_150_0(core__GEN_150_0),
    ._GEN_283(core__GEN_283),
    ._GEN_184(core__GEN_184),
    ._GEN_178_0(core__GEN_178_0),
    ._GEN_68_0(core__GEN_68_0),
    ._GEN_296_0(core__GEN_296_0),
    ._GEN_382(core__GEN_382),
    ._GEN_397(core__GEN_397),
    ._GEN_277(core__GEN_277),
    ._GEN_395_0(core__GEN_395_0),
    ._GEN_304_0(core__GEN_304_0),
    ._GEN_199(core__GEN_199),
    ._GEN_403(core__GEN_403),
    ._GEN_262(core__GEN_262),
    ._GEN_28(core__GEN_28),
    ._GEN_275_0(core__GEN_275_0),
    ._GEN_269_0(core__GEN_269_0),
    ._GEN_361(core__GEN_361),
    ._GEN_96(core__GEN_96),
    ._GEN_278_0(core__GEN_278_0),
    ._GEN_193(core__GEN_193),
    ._GEN_379(core__GEN_379),
    ._GEN_244_0(core__GEN_244_0),
    ._GEN_138(core__GEN_138),
    ._GEN_271(core__GEN_271),
    ._GEN_251_0(core__GEN_251_0),
    ._GEN_151_1(core__GEN_151_1),
    ._GEN_166_0(core__GEN_166_0),
    ._GEN_455(core__GEN_455),
    ._GEN_370(core__GEN_370),
    ._GEN_364(core__GEN_364),
    ._GEN_259(core__GEN_259),
    ._GEN_377_0(core__GEN_377_0),
    ._GEN_153_0(core__GEN_153_0),
    ._GEN_292(core__GEN_292),
    ._GEN_84(core__GEN_84),
    ._GEN_78(core__GEN_78),
    ._GEN_272_0(core__GEN_272_0),
    ._GEN_47_0(core__GEN_47_0),
    ._GEN_335_0(core__GEN_335_0),
    ._GEN_41_0(core__GEN_41_0),
    ._GEN_385(core__GEN_385),
    ._GEN_250(core__GEN_250),
    ._GEN_434(core__GEN_434),
    ._GEN_257_0(core__GEN_257_0),
    ._GEN_343(core__GEN_343),
    ._GEN_443(core__GEN_443),
    ._GEN_105(core__GEN_105),
    ._GEN_99(core__GEN_99),
    ._GEN_358(core__GEN_358),
    ._GEN_356_0(core__GEN_356_0),
    ._GEN_350_0(core__GEN_350_0),
    ._GEN_132_0(core__GEN_132_0),
    ._GEN_22(core__GEN_22),
    ._GEN_144(core__GEN_144),
    ._GEN_265(core__GEN_265),
    ._GEN_17(core__GEN_17),
    ._GEN_159(core__GEN_159),
    ._GEN_428(core__GEN_428),
    ._GEN_449(core__GEN_449),
    ._GEN_90_0(core__GEN_90_0),
    ._GEN_172_0(core__GEN_172_0),
    ._GEN_187(core__GEN_187),
    ._GEN_117_0(core__GEN_117_0),
    ._GEN_236_0(core__GEN_236_0),
    ._GEN_371_0(core__GEN_371_0),
    ._GEN_391(core__GEN_391),
    ._GEN_165(core__GEN_165),
    ._GEN_286(core__GEN_286),
    ._GEN_145_0(core__GEN_145_0),
    ._GEN_284_0(core__GEN_284_0),
    ._GEN_232(core__GEN_232),
    ._GEN_147_0(core__GEN_147_0),
    ._GEN_416_0(core__GEN_416_0),
    ._GEN_274(core__GEN_274),
    ._GEN_260_0(core__GEN_260_0),
    ._GEN_175_0(core__GEN_175_0),
    ._GEN_105_0(core__GEN_105_0),
    ._GEN_169_0(core__GEN_169_0),
    ._GEN_338_0(core__GEN_338_0),
    ._GEN_247(core__GEN_247),
    ._GEN_133_0(core__GEN_133_0),
    ._GEN_141_0(core__GEN_141_0),
    ._GEN_160_0(core__GEN_160_0),
    ._GEN_346(core__GEN_346),
    ._GEN_99_0(core__GEN_99_0),
    ._GEN_344_0(core__GEN_344_0),
    ._GEN_373(core__GEN_373),
    ._GEN_424_0(core__GEN_424_0),
    ._GEN_239_0(core__GEN_239_0),
    ._GEN_353_0(core__GEN_353_0),
    ._GEN_268(core__GEN_268),
    ._GEN_127_0(core__GEN_127_0),
    ._GEN_8(core__GEN_8),
    ._GEN_266_0(core__GEN_266_0),
    ._GEN_331_0(core__GEN_331_0),
    ._GEN_452(core__GEN_452),
    ._GEN_93_0(core__GEN_93_0),
    ._GEN_87_0(core__GEN_87_0),
    ._GEN_367(core__GEN_367),
    ._GEN_226(core__GEN_226),
    ._GEN_120_0(core__GEN_120_0),
    ._GEN_365_0(core__GEN_365_0),
    ._GEN_6(core__GEN_6),
    ._GEN_410_0(core__GEN_410_0),
    ._GEN_253_0(core__GEN_253_0),
    ._GEN_152_0(core__GEN_152_0),
    ._GEN_325_0(core__GEN_325_0),
    ._GEN_148_0(core__GEN_148_0),
    ._GEN_437(core__GEN_437),
    ._GEN_352_0(core__GEN_352_0),
    ._GEN_332_0(core__GEN_332_0),
    ._GEN_108(core__GEN_108),
    ._GEN_126_0(core__GEN_126_0),
    ._GEN_245_0(core__GEN_245_0),
    ._GEN_359_0(core__GEN_359_0),
    ._GEN_431(core__GEN_431),
    ._GEN_72_0(core__GEN_72_0),
    ._GEN_66(core__GEN_66),
    ._GEN_154_0(core__GEN_154_0),
    ._GEN_458(core__GEN_458),
    ._GEN_317_0(core__GEN_317_0),
    ._GEN_326_0(core__GEN_326_0),
    ._GEN_241(core__GEN_241),
    ._GEN_341_0(core__GEN_341_0),
    ._GEN_402_0(core__GEN_402_0),
    ._GEN_1_2(core__GEN_1_2),
    ._GEN_48(core__GEN_48),
    ._GEN_394_0(core__GEN_394_0),
    ._GEN_60(core__GEN_60),
    ._GEN_248_0(core__GEN_248_0),
    ._GEN_75_0(core__GEN_75_0),
    ._GEN_349(core__GEN_349),
    ._GEN_214(core__GEN_214),
    ._GEN_347_0(core__GEN_347_0),
    ._GEN_412_0(core__GEN_412_0),
    ._GEN_92_0(core__GEN_92_0),
    ._GEN_102_0(core__GEN_102_0),
    ._GEN_256(core__GEN_256),
    ._GEN_121_0(core__GEN_121_0),
    ._GEN_425_0(core__GEN_425_0),
    ._GEN_305_0(core__GEN_305_0),
    ._GEN_419_0(core__GEN_419_0),
    ._GEN_81(core__GEN_81),
    ._GEN_320_0(core__GEN_320_0),
    ._GEN_108_0(core__GEN_108_0),
    ._GEN_114_0(core__GEN_114_0),
    ._GEN_123_0(core__GEN_123_0),
    ._GEN_413_0(core__GEN_413_0),
    ._GEN_54(core__GEN_54),
    ._GEN_136_0(core__GEN_136_0),
    ._GEN_142_0(core__GEN_142_0),
    ._GEN_440(core__GEN_440),
    ._GEN_295_0(core__GEN_295_0),
    ._GEN_340(core__GEN_340),
    ._GEN_355(core__GEN_355),
    ._GEN_235(core__GEN_235),
    ._GEN_129_0(core__GEN_129_0),
    ._GEN_404_0(core__GEN_404_0),
    ._GEN_403_0(core__GEN_403_0),
    ._GEN_313_0(core__GEN_313_0),
    ._GEN_242_0(core__GEN_242_0),
    ._GEN_69_0(core__GEN_69_0),
    ._GEN_157_0(core__GEN_157_0),
    ._GEN_220(core__GEN_220),
    ._GEN_229(core__GEN_229),
    ._GEN_115_0(core__GEN_115_0),
    ._GEN_15_0(core__GEN_15_0),
    ._GEN_334(core__GEN_334),
    ._GEN_328(core__GEN_328),
    ._GEN_96_0(core__GEN_96_0),
    ._GEN_86_0(core__GEN_86_0),
    ._GEN_36(core__GEN_36),
    ._GEN_405_0(core__GEN_405_0),
    ._GEN_415_0(core__GEN_415_0),
    ._GEN_164_0(core__GEN_164_0),
    ._GEN_124_0(core__GEN_124_0),
    ._GEN_322(core__GEN_322),
    ._GEN_308_0(core__GEN_308_0),
    ._GEN_337_0(core__GEN_337_0),
    ._GEN_223(core__GEN_223),
    ._GEN_217(core__GEN_217),
    ._GEN_192(core__GEN_192),
    ._GEN_390_0(core__GEN_390_0),
    ._GEN_42_0(core__GEN_42_0),
    ._GEN_149_0(core__GEN_149_0),
    ._GEN_291_0(core__GEN_291_0),
    ._GEN_139_0(core__GEN_139_0),
    ._GEN_329_0(core__GEN_329_0),
    ._GEN_292_0(core__GEN_292_0),
    ._GEN_298_0(core__GEN_298_0),
    ._GEN_207(core__GEN_207),
    ._GEN_399_0(core__GEN_399_0),
    ._GEN_421(core__GEN_421),
    ._GEN_63(core__GEN_63),
    ._GEN_391_0(core__GEN_391_0),
    ._GEN_316_0(core__GEN_316_0),
    ._GEN_306_0(core__GEN_306_0),
    ._GEN_314_0(core__GEN_314_0),
    ._GEN_21_0(core__GEN_21_0),
    ._GEN_323_0(core__GEN_323_0),
    ._GEN_384_0(core__GEN_384_0),
    ._GEN_118_0(core__GEN_118_0),
    ._GEN_376_0(core__GEN_376_0),
    ._GEN_422_0(core__GEN_422_0),
    ._GEN_277_0(core__GEN_277_0),
    ._GEN_57(core__GEN_57),
    ._GEN_130_0(core__GEN_130_0),
    ._GEN_46_0(core__GEN_46_0),
    ._GEN_111_0(core__GEN_111_0),
    ._GEN_78_0(core__GEN_78_0),
    ._GEN_238_0(core__GEN_238_0),
    ._GEN_407_0(core__GEN_407_0),
    ._GEN_179_0(core__GEN_179_0),
    ._GEN_397_0(core__GEN_397_0),
    ._GEN_173_0(core__GEN_173_0),
    ._GEN_70_0(core__GEN_70_0),
    ._GEN_379_0(core__GEN_379_0),
    ._GEN_82_0(core__GEN_82_0),
    ._GEN_373_0(core__GEN_373_0),
    ._GEN_45_0(core__GEN_45_0),
    ._GEN_54_0(core__GEN_54_0),
    ._GEN_201(core__GEN_201),
    ._GEN_195(core__GEN_195),
    ._GEN_364_0(core__GEN_364_0),
    ._GEN_259_0(core__GEN_259_0),
    ._GEN_167_0(core__GEN_167_0),
    ._GEN_309_0(core__GEN_309_0),
    ._GEN_43_0(core__GEN_43_0),
    ._GEN_372_0(core__GEN_372_0),
    ._GEN_19(core__GEN_19),
    ._GEN_161_0(core__GEN_161_0),
    ._GEN_51(core__GEN_51),
    ._GEN_265_0(core__GEN_265_0),
    ._GEN_294_0(core__GEN_294_0),
    ._GEN_180(core__GEN_180),
    ._GEN_189(core__GEN_189),
    ._GEN_211(core__GEN_211),
    ._GEN_301_0(core__GEN_301_0),
    ._GEN_393_0(core__GEN_393_0),
    ._GEN_387_0(core__GEN_387_0),
    ._GEN_39(core__GEN_39),
    ._GEN_146_1(core__GEN_146_1),
    ._GEN_288_0(core__GEN_288_0),
    ._GEN_310_0(core__GEN_310_0),
    ._GEN_300_0(core__GEN_300_0),
    ._GEN_286_0(core__GEN_286_0),
    ._GEN_400_0(core__GEN_400_0),
    ._GEN_319_0(core__GEN_319_0),
    ._GEN_107_0(core__GEN_107_0),
    ._GEN_174_0(core__GEN_174_0),
    ._GEN_89(core__GEN_89),
    ._GEN_358_0(core__GEN_358_0),
    ._GEN_30(core__GEN_30),
    ._GEN_24(core__GEN_24),
    ._GEN_408_0(core__GEN_408_0),
    ._GEN_418_0(core__GEN_418_0),
    ._GEN_273_0(core__GEN_273_0),
    ._GEN_5_0(core__GEN_5_0),
    ._GEN_112_0(core__GEN_112_0),
    ._GEN_385_0(core__GEN_385_0),
    ._GEN_457(core__GEN_457),
    ._GEN_311_0(core__GEN_311_0),
    ._GEN_280_0(core__GEN_280_0),
    ._GEN_366_0(core__GEN_366_0),
    ._GEN_360_0(core__GEN_360_0),
    ._GEN_354_0(core__GEN_354_0),
    ._GEN_143_0(core__GEN_143_0),
    ._GEN_367_0(core__GEN_367_0),
    ._GEN_33_0(core__GEN_33_0),
    ._GEN_247_0(core__GEN_247_0),
    ._GEN_276_0(core__GEN_276_0),
    ._GEN_348_0(core__GEN_348_0),
    ._GEN_274_0(core__GEN_274_0),
    ._GEN_460(core__GEN_460),
    ._GEN_101_0(core__GEN_101_0),
    ._GEN_375_0(core__GEN_375_0),
    ._GEN_283_0(core__GEN_283_0),
    ._GEN_27(core__GEN_27),
    ._GEN_13(core__GEN_13),
    ._GEN_388_0(core__GEN_388_0),
    ._GEN_382_0(core__GEN_382_0),
    ._GEN_268_0(core__GEN_268_0),
    ._GEN_297_0(core__GEN_297_0),
    ._GEN_89_0(core__GEN_89_0),
    ._GEN_176_0(core__GEN_176_0),
    ._GEN_177_0(core__GEN_177_0),
    ._GEN_346_0(core__GEN_346_0),
    ._GEN_64_0(core__GEN_64_0),
    ._GEN_340_0(core__GEN_340_0),
    ._GEN_255_0(core__GEN_255_0),
    ._GEN_204(core__GEN_204),
    ._GEN_134_0(core__GEN_134_0),
    ._GEN_149_1(core__GEN_149_1),
    ._GEN_439(core__GEN_439),
    ._GEN_80_0(core__GEN_80_0),
    ._GEN_262_0(core__GEN_262_0),
    ._GEN_303_0(core__GEN_303_0),
    ._GEN_162_0(core__GEN_162_0),
    ._GEN_17_0(core__GEN_17_0),
    ._GEN_198(core__GEN_198),
    ._GEN_361_0(core__GEN_361_0),
    ._GEN_381_0(core__GEN_381_0),
    ._GEN_261_0(core__GEN_261_0),
    ._GEN_155_0(core__GEN_155_0),
    ._GEN_156_0(core__GEN_156_0),
    ._GEN_170_0(core__GEN_170_0),
    ._GEN_95_0(core__GEN_95_0),
    ._GEN_183(core__GEN_183),
    ._GEN_369_0(core__GEN_369_0),
    ._GEN_73_0(core__GEN_73_0),
    ._GEN_128_0(core__GEN_128_0),
    ._GEN_241_0(core__GEN_241_0),
    ._GEN_282_0(core__GEN_282_0),
    ._GEN_396_0(core__GEN_396_0),
    ._GEN_445(core__GEN_445),
    ._GEN_289_0(core__GEN_289_0),
    ._GEN_378_0(core__GEN_378_0),
    ._GEN_186(core__GEN_186),
    ._GEN_131_0(core__GEN_131_0),
    ._GEN_152_1(core__GEN_152_1),
    ._GEN_421_0(core__GEN_421_0),
    ._GEN_427(core__GEN_427),
    ._GEN_62(core__GEN_62),
    ._GEN_285_0(core__GEN_285_0),
    ._GEN_336_0(core__GEN_336_0),
    ._GEN_144_0(core__GEN_144_0),
    ._GEN_150_1(core__GEN_150_1),
    ._GEN_454(core__GEN_454),
    ._GEN_363_0(core__GEN_363_0),
    ._GEN_243_0(core__GEN_243_0),
    ._GEN_258_0(core__GEN_258_0),
    ._GEN_138_0(core__GEN_138_0),
    ._GEN_256_0(core__GEN_256_0),
    ._GEN_171_0(core__GEN_171_0),
    ._GEN_357_0(core__GEN_357_0),
    ._GEN_165_0(core__GEN_165_0),
    ._GEN_110_0(core__GEN_110_0),
    ._GEN_40_0(core__GEN_40_0),
    ._GEN_264_0(core__GEN_264_0),
    ._GEN_5_1(core__GEN_5_1),
    ._GEN_158_0(core__GEN_158_0),
    ._GEN_16_0(core__GEN_16_0),
    ._GEN_271_0(core__GEN_271_0),
    ._GEN_342_0(core__GEN_342_0),
    ._GEN_322_0(core__GEN_322_0),
    ._GEN_98_0(core__GEN_98_0),
    ._GEN_237_0(core__GEN_237_0),
    ._GEN_334_0(core__GEN_334_0),
    ._GEN_116_0(core__GEN_116_0),
    ._GEN_235_0(core__GEN_235_0),
    ._GEN_349_0(core__GEN_349_0),
    ._GEN_147_1(core__GEN_147_1),
    ._GEN_448(core__GEN_448),
    ._GEN_442(core__GEN_442),
    ._GEN_83_0(core__GEN_83_0),
    ._GEN_343_0(core__GEN_343_0),
    ._GEN_355_0(core__GEN_355_0),
    ._GEN_137_0(core__GEN_137_0),
    ._GEN_370_0(core__GEN_370_0),
    ._GEN_250_0(core__GEN_250_0),
    ._GEN_77(core__GEN_77),
    ._GEN_270_0(core__GEN_270_0),
    ._GEN_279_0(core__GEN_279_0),
    ._GEN_159_0(core__GEN_159_0),
    ._GEN_463(core__GEN_463),
    ._GEN_328_0(core__GEN_328_0),
    ._GEN_104_0(core__GEN_104_0)
  );
  AsyncScratchPadMemory memory ( // @[top.scala 24:28]
    .metaReset(memory_metaReset),
    .clock(memory_clock),
    .io_core_ports_0_req_valid(memory_io_core_ports_0_req_valid),
    .io_core_ports_0_req_bits_addr(memory_io_core_ports_0_req_bits_addr),
    .io_core_ports_0_req_bits_data(memory_io_core_ports_0_req_bits_data),
    .io_core_ports_0_req_bits_fcn(memory_io_core_ports_0_req_bits_fcn),
    .io_core_ports_0_req_bits_typ(memory_io_core_ports_0_req_bits_typ),
    .io_core_ports_0_resp_valid(memory_io_core_ports_0_resp_valid),
    .io_core_ports_0_resp_bits_data(memory_io_core_ports_0_resp_bits_data),
    ._GEN_4_0(memory__GEN_4_0),
    ._GEN_1_1(memory__GEN_1_1),
    ._GEN_0_1(memory__GEN_0_1),
    ._GEN_3_1(memory__GEN_3_1),
    ._GEN_5_0(memory__GEN_5_0),
    ._GEN_2_0(memory__GEN_2_0)
  );
  assign core_metaReset = metaReset;
  assign memory_metaReset = metaReset;
  assign io_imem_req_valid = 1'h1; // @[top.scala 29:22]
  assign io_imem_req_bits_addr = core_io_imem_req_bits_addr; // @[top.scala 29:22]
  assign io_imem_req_bits_data = 32'h0; // @[top.scala 29:22]
  assign io_imem_req_bits_fcn = 1'h0; // @[top.scala 29:22]
  assign io_imem_req_bits_typ = 3'h0; // @[top.scala 29:22]
  assign assert_out = core__GEN_463;
  assign auto_cover_out = {_GEN_1584,profilePin_791};
  assign core_clock = clock;
  assign core_reset = reset; // @[top.scala 35:20]
  assign core_io_imem_resp_valid = io_imem_resp_valid; // @[top.scala 29:22]
  assign core_io_imem_resp_bits_data = io_imem_resp_bits_data; // @[top.scala 29:22]
  assign core_io_dmem_resp_valid = memory_io_core_ports_0_resp_valid; // @[top.scala 28:22]
  assign core_io_dmem_resp_bits_data = memory_io_core_ports_0_resp_bits_data; // @[top.scala 28:22]
  assign memory_clock = clock;
  assign memory_io_core_ports_0_req_valid = core_io_dmem_req_valid; // @[top.scala 28:22]
  assign memory_io_core_ports_0_req_bits_addr = core_io_dmem_req_bits_addr; // @[top.scala 28:22]
  assign memory_io_core_ports_0_req_bits_data = core_io_dmem_req_bits_data; // @[top.scala 28:22]
  assign memory_io_core_ports_0_req_bits_fcn = core_io_dmem_req_bits_fcn; // @[top.scala 28:22]
  assign memory_io_core_ports_0_req_bits_typ = core_io_dmem_req_bits_typ; // @[top.scala 28:22]
endmodule
module CtlPath(
  input         metaReset,
  input         clock,
  input         reset,
  input         io_imem_resp_valid,
  input         io_dmem_resp_valid,
  input  [31:0] io_dat_dec_inst,
  input         io_dat_exe_br_eq,
  input         io_dat_exe_br_lt,
  input         io_dat_exe_br_ltu,
  input  [3:0]  io_dat_exe_br_type,
  input         io_dat_mem_ctrl_dmem_val,
  input         io_dat_csr_eret,
  output        io_ctl_dec_stall,
  output        io_ctl_full_stall,
  output [1:0]  io_ctl_exe_pc_sel,
  output [3:0]  io_ctl_br_type,
  output        io_ctl_if_kill,
  output        io_ctl_dec_kill,
  output [1:0]  io_ctl_op1_sel,
  output [2:0]  io_ctl_op2_sel,
  output [3:0]  io_ctl_alu_fun,
  output [1:0]  io_ctl_wb_sel,
  output        io_ctl_rf_wen,
  output        io_ctl_mem_val,
  output [1:0]  io_ctl_mem_fcn,
  output [2:0]  io_ctl_mem_typ,
  output [2:0]  io_ctl_csr_cmd,
  output        io_ctl_fencei,
  output        io_ctl_pipeline_kill,
  output        io_ctl_mem_exception,
  output        _GEN_111_0,
  output        _GEN_71_0,
  output        _GEN_324_0,
  output        _GEN_219_0,
  output        _GEN_168_0,
  output        _GEN_1_0,
  output        _GEN_423_0,
  output        _GEN_44_0,
  output        _GEN_267_0,
  output        _GEN_126_0,
  output        _GEN_153_0,
  output        _GEN_225_0,
  output        _GEN_59_0,
  output        _GEN_252_0,
  output        _GEN_147_0,
  output        _GEN_351_0,
  output        _GEN_210_0,
  output        _GEN_246_0,
  output        _GEN_65_0,
  output        _GEN_132_0,
  output        _GEN_318_0,
  output        _GEN_92_0,
  output        _GEN_345_0,
  output        _GEN_231_0,
  output        _GEN_417_0,
  output        _GEN_50_0,
  output        _GEN_330_0,
  output        _GEN_86_0,
  output        _GEN_339_0,
  output        _GEN_240_0,
  output        _GEN_234_0,
  output        _GEN_120_0,
  output        _GEN_129_0,
  output        _GEN_333_0,
  output        _GEN_302_0,
  output        _GEN_228_0,
  output        _GEN_197_0,
  output        _GEN_411_0,
  output        _GEN_401_0,
  output        _GEN_47_0,
  output        _GEN_296_0,
  output        _GEN_74_0,
  output        _GEN_213_0,
  output        _GEN_32_0,
  output        _GEN_68_0,
  output        _GEN_135_0,
  output        _GEN_26_0,
  output        _GEN_53_0,
  output        _GEN_141_0,
  output        _GEN_327_0,
  output        _GEN_395_0,
  output        _GEN_249_0,
  output        _GEN_114_0,
  output        _GEN_312_0,
  output        _GEN_203_0,
  output        _GEN_20_0,
  output        _GEN_15_0,
  output        _GEN_216_0,
  output        _GEN_206_0,
  output        _GEN_420_0,
  output        _GEN_123_0,
  output        _GEN_315_0,
  output        _GEN_284_0,
  output        _GEN_179_0,
  output        _GEN_222_0,
  output        _GEN_377_0,
  output        _GEN_191_0,
  output        _GEN_290_0,
  output        _GEN_404_0,
  output        _GEN_56_1,
  output        _GEN_305_0,
  output        _GEN_299_0,
  output        _GEN_185_0,
  output        _GEN_398_0,
  output        _GEN_41_0,
  output        _GEN_321_0,
  output        _GEN_414_0,
  output        _GEN_383_0,
  output        _GEN_35_0,
  output        _GEN_29_0,
  output        _GEN_278_0,
  output        _GEN_117_0,
  output        _GEN_365_0,
  output        _GEN_359_0,
  output        _GEN_38_0,
  output        _GEN_167_0,
  output        _GEN_350_0,
  output        _GEN_106_0,
  output        _GEN_18_0,
  output        _GEN_293_0,
  output        _GEN_371_0,
  output        _GEN_251_0,
  output        _GEN_209_0,
  output        _GEN_308_0,
  output        _GEN_173_0,
  output        _GEN_200_0,
  output        _GEN_386_0,
  output        _GEN_272_0,
  output        _GEN_91_1,
  output        _GEN_194_0,
  output        _GEN_188_0,
  output        _GEN_392_0,
  output        _GEN_23_0,
  output        _GEN_407_0,
  output        _GEN_287_0,
  output        _GEN_266_0,
  output        _GEN_374_0,
  output        _GEN_233_0,
  output        _GEN_269_0,
  output        _GEN_260_0,
  output        _GEN_161_0,
  output        _GEN_155_0,
  output        _GEN_368_0,
  output        _GEN_254_0,
  output        _GEN_281_0,
  output        _GEN_73_0,
  output        _GEN_353_0,
  output        _GEN_332_0,
  output        _GEN_88_1,
  output        _GEN_176_0,
  output        _GEN_380_0,
  output        _GEN_389_0,
  output        _GEN_94_0,
  output        _GEN_347_0,
  output        _GEN_109_0,
  output        _GEN_182_0,
  output        _GEN_9_0,
  output        _GEN_149_0,
  output        _GEN_248_0,
  output        _GEN_275_0,
  output        _GEN_140_1,
  output        _GEN_100_0,
  output        _GEN_362_0,
  output        _GEN_413_0,
  output        _GEN_76_0,
  output        _GEN_164_0,
  output        _GEN_242_0,
  output        _GEN_137_0,
  output        _GEN_341_0,
  output        _GEN_263_0,
  output        _GEN_257_0,
  output        _GEN_122_1,
  output        _GEN_143_0,
  output        _GEN_82_0,
  output        _GEN_170_0,
  output        _GEN_356_0,
  output        _GEN_221_0,
  output        _GEN_215_0,
  output        _GEN_320_0,
  output        _GEN_314_0,
  output        _GEN_329_0,
  output        _GEN_103_1,
  output        _GEN_97_0,
  output        _GEN_236_0,
  output        _GEN_61_0,
  output        _GEN_55_0,
  output        _GEN_335_0,
  output        _GEN_158_0,
  output        _GEN_422_0,
  output        _GEN_245_0,
  output        _GEN_37_0,
  output        _GEN_125_1,
  output        _GEN_70_0,
  output        _GEN_64_0,
  output        _GEN_344_0,
  output        _GEN_338_0,
  output        _GEN_416_0,
  output        _GEN_406_1,
  output        _GEN_58_0,
  output        _GEN_85_1,
  output        _GEN_43_0,
  output        _GEN_131_0,
  output        _GEN_230_0,
  output        _GEN_239_0,
  output        _GEN_152_0,
  output        _GEN_307_1,
  output        _GEN_146_1,
  output        _GEN_224_0,
  output        _GEN_110_0,
  output        _GEN_119_1,
  output        _GEN_323_0,
  output        _GEN_317_0,
  output        _GEN_79_1,
  output        _GEN_218_0,
  output        _GEN_208_0,
  output        _GEN_196_0,
  output        _GEN_31_0,
  output        _GEN_400_0,
  output        _GEN_113_1,
  output        _GEN_212_0,
  output        _GEN_181_0,
  output        _GEN_227_0,
  output        _GEN_425_0,
  output        _GEN_280_0,
  output        _GEN_46_0,
  output        _GEN_134_0,
  output        _GEN_289_0,
  output        _GEN_202_0,
  output        _GEN_419_0,
  output        _GEN_388_0,
  output        _GEN_410_0,
  output        _GEN_52_0,
  output        _GEN_311_0,
  output        _GEN_301_0,
  output        _GEN_295_0,
  output        _GEN_67_0,
  output        _GEN_25_0,
  output        _GEN_409_1,
  output        _GEN_326_0,
  output        _GEN_394_0,
  output        _GEN_128_0,
  output        _GEN_376_0,
  output        _GEN_40_0,
  output        _GEN_34_0,
  output        _GEN_49_0,
  output        _GEN_102_0,
  output        _GEN_190_0,
  output        _GEN_205_0,
  output        _GEN_298_0,
  output        _GEN_163_1,
  output        _GEN_14_0,
  output        _GEN_116_0,
  output        _GEN_283_0,
  output        _GEN_184_0,
  output        _GEN_178_1,
  output        _GEN_382_0,
  output        _GEN_397_0,
  output        _GEN_277_0,
  output        _GEN_304_1,
  output        _GEN_199_0,
  output        _GEN_403_0,
  output        _GEN_262_0,
  output        _GEN_28_0,
  output        _GEN_361_0,
  output        _GEN_96_0,
  output        _GEN_193_0,
  output        _GEN_379_0,
  output        _GEN_244_1,
  output        _GEN_271_0,
  output        _GEN_151_2,
  output        _GEN_166_1,
  output        _GEN_370_0,
  output        _GEN_364_0,
  output        _GEN_259_0,
  output        _GEN_292_0,
  output        _GEN_84_0,
  output        _GEN_78_0,
  output        _GEN_385_0,
  output        _GEN_250_0,
  output        _GEN_343_0,
  output        _GEN_105_0,
  output        _GEN_99_0,
  output        _GEN_358_0,
  output        _GEN_22_0,
  output        _GEN_265_0,
  output        _GEN_17_0,
  output        _GEN_90_1,
  output        _GEN_172_1,
  output        _GEN_187_0,
  output        _GEN_391_0,
  output        _GEN_286_0,
  output        _GEN_145_1,
  output        _GEN_232_0,
  output        _GEN_274_0,
  output        _GEN_175_1,
  output        _GEN_169_1,
  output        _GEN_247_0,
  output        _GEN_133_1,
  output        _GEN_160_1,
  output        _GEN_346_0,
  output        _GEN_373_0,
  output        _GEN_424_1,
  output        _GEN_268_0,
  output        _GEN_127_1,
  output        _GEN_8_0,
  output        _GEN_331_1,
  output        _GEN_93_1,
  output        _GEN_87_1,
  output        _GEN_367_0,
  output        _GEN_226_0,
  output        _GEN_253_1,
  output        _GEN_325_1,
  output        _GEN_148_1,
  output        _GEN_352_1,
  output        _GEN_108_0,
  output        _GEN_72_1,
  output        _GEN_66_0,
  output        _GEN_154_1,
  output        _GEN_241_0,
  output        _GEN_402_1,
  output        _GEN_48_0,
  output        _GEN_60_0,
  output        _GEN_75_1,
  output        _GEN_349_0,
  output        _GEN_214_0,
  output        _GEN_412_1,
  output        _GEN_256_0,
  output        _GEN_121_1,
  output        _GEN_81_0,
  output        _GEN_54_0,
  output        _GEN_136_1,
  output        _GEN_142_1,
  output        _GEN_340_0,
  output        _GEN_355_0,
  output        _GEN_235_0,
  output        _GEN_313_1,
  output        _GEN_69_1,
  output        _GEN_157_1,
  output        _GEN_220_0,
  output        _GEN_229_0,
  output        _GEN_115_1,
  output        _GEN_334_0,
  output        _GEN_328_0,
  output        _GEN_36_0,
  output        _GEN_405_1,
  output        _GEN_415_1,
  output        _GEN_124_1,
  output        _GEN_322_0,
  output        _GEN_337_1,
  output        _GEN_223_0,
  output        _GEN_217_0,
  output        _GEN_192_0,
  output        _GEN_390_1,
  output        _GEN_42_1,
  output        _GEN_291_1,
  output        _GEN_139_1,
  output        _GEN_207_0,
  output        _GEN_399_1,
  output        _GEN_421_0,
  output        _GEN_63_0,
  output        _GEN_316_1,
  output        _GEN_306_1,
  output        _GEN_21_1,
  output        _GEN_384_1,
  output        _GEN_118_1,
  output        _GEN_57_0,
  output        _GEN_130_1,
  output        _GEN_238_1,
  output        _GEN_45_1,
  output        _GEN_201_0,
  output        _GEN_195_0,
  output        _GEN_309_1,
  output        _GEN_372_1,
  output        _GEN_19_0,
  output        _GEN_51_0,
  output        _GEN_294_1,
  output        _GEN_180_0,
  output        _GEN_189_0,
  output        _GEN_211_0,
  output        _GEN_393_1,
  output        _GEN_387_1,
  output        _GEN_39_0,
  output        _GEN_288_1,
  output        _GEN_310_1,
  output        _GEN_300_1,
  output        _GEN_319_1,
  output        _GEN_107_1,
  output        _GEN_174_1,
  output        _GEN_30_0,
  output        _GEN_24_0,
  output        _GEN_408_1,
  output        _GEN_418_1,
  output        _GEN_273_1,
  output        _GEN_5_1,
  output        _GEN_112_1,
  output        _GEN_366_1,
  output        _GEN_360_1,
  output        _GEN_354_1,
  output        _GEN_33_1,
  output        _GEN_276_1,
  output        _GEN_348_1,
  output        _GEN_101_1,
  output        _GEN_375_1,
  output        _GEN_27_0,
  output        _GEN_13_0,
  output        _GEN_297_1,
  output        _GEN_89_1,
  output        _GEN_177_1,
  output        _GEN_255_1,
  output        _GEN_204_0,
  output        _GEN_80_1,
  output        _GEN_303_1,
  output        _GEN_162_1,
  output        _GEN_198_0,
  output        _GEN_381_1,
  output        _GEN_261_1,
  output        _GEN_156_1,
  output        _GEN_95_1,
  output        _GEN_183_0,
  output        _GEN_369_1,
  output        _GEN_282_1,
  output        _GEN_396_1,
  output        _GEN_378_1,
  output        _GEN_186_0,
  output        _GEN_62_0,
  output        _GEN_285_1,
  output        _GEN_336_1,
  output        _GEN_144_1,
  output        _GEN_150_2,
  output        _GEN_363_1,
  output        _GEN_243_1,
  output        _GEN_258_1,
  output        _GEN_138_1,
  output        _GEN_171_1,
  output        _GEN_357_1,
  output        _GEN_165_1,
  output        _GEN_264_1,
  output        _GEN_16_1,
  output        _GEN_342_1,
  output        _GEN_98_1,
  output        _GEN_237_1,
  output        _GEN_83_1,
  output        _GEN_77_0,
  output        _GEN_270_1,
  output        _GEN_279_1,
  output        _GEN_159_1,
  output        _GEN_104_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] _T_232 = io_dat_dec_inst & 32'h707f; // @[Lookup.scala 9:38]
  wire  _T_233 = 32'h2003 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_237 = 32'h3 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_241 = 32'h4003 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_245 = 32'h1003 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_249 = 32'h5003 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_253 = 32'h2023 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_257 = 32'h23 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_261 = 32'h1023 == _T_232; // @[Lookup.scala 9:38]
  wire [31:0] _T_264 = io_dat_dec_inst & 32'h7f; // @[Lookup.scala 9:38]
  wire  _T_265 = 32'h17 == _T_264; // @[Lookup.scala 9:38]
  wire  _T_269 = 32'h37 == _T_264; // @[Lookup.scala 9:38]
  wire  _T_273 = 32'h13 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_277 = 32'h7013 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_281 = 32'h6013 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_285 = 32'h4013 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_289 = 32'h2013 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_293 = 32'h3013 == _T_232; // @[Lookup.scala 9:38]
  wire [31:0] _T_296 = io_dat_dec_inst & 32'hfc00707f; // @[Lookup.scala 9:38]
  wire  _T_297 = 32'h1013 == _T_296; // @[Lookup.scala 9:38]
  wire  _T_301 = 32'h40005013 == _T_296; // @[Lookup.scala 9:38]
  wire  _T_305 = 32'h5013 == _T_296; // @[Lookup.scala 9:38]
  wire [31:0] _T_308 = io_dat_dec_inst & 32'hfe00707f; // @[Lookup.scala 9:38]
  wire  _T_309 = 32'h1033 == _T_308; // @[Lookup.scala 9:38]
  wire  _T_313 = 32'h33 == _T_308; // @[Lookup.scala 9:38]
  wire  _T_317 = 32'h40000033 == _T_308; // @[Lookup.scala 9:38]
  wire  _T_321 = 32'h2033 == _T_308; // @[Lookup.scala 9:38]
  wire  _T_325 = 32'h3033 == _T_308; // @[Lookup.scala 9:38]
  wire  _T_329 = 32'h7033 == _T_308; // @[Lookup.scala 9:38]
  wire  _T_333 = 32'h6033 == _T_308; // @[Lookup.scala 9:38]
  wire  _T_337 = 32'h4033 == _T_308; // @[Lookup.scala 9:38]
  wire  _T_341 = 32'h40005033 == _T_308; // @[Lookup.scala 9:38]
  wire  _T_345 = 32'h5033 == _T_308; // @[Lookup.scala 9:38]
  wire  _T_349 = 32'h6f == _T_264; // @[Lookup.scala 9:38]
  wire  _T_353 = 32'h67 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_357 = 32'h63 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_361 = 32'h1063 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_365 = 32'h5063 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_369 = 32'h7063 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_373 = 32'h4063 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_377 = 32'h6063 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_381 = 32'h5073 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_385 = 32'h6073 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_389 = 32'h1073 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_393 = 32'h2073 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_397 = 32'h3073 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_401 = 32'h7073 == _T_232; // @[Lookup.scala 9:38]
  wire  _T_405 = 32'h73 == io_dat_dec_inst; // @[Lookup.scala 9:38]
  wire  _T_409 = 32'h30200073 == io_dat_dec_inst; // @[Lookup.scala 9:38]
  wire  _T_413 = 32'h7b200073 == io_dat_dec_inst; // @[Lookup.scala 9:38]
  wire  _T_417 = 32'h100073 == io_dat_dec_inst; // @[Lookup.scala 9:38]
  wire  _T_421 = 32'h10500073 == io_dat_dec_inst; // @[Lookup.scala 9:38]
  wire  _T_425 = 32'h100f == _T_232; // @[Lookup.scala 9:38]
  wire  _T_429 = 32'hf == _T_232; // @[Lookup.scala 9:38]
  wire  _T_431 = _T_425 | _T_429; // @[Lookup.scala 11:37]
  wire  _T_432 = _T_421 | _T_431; // @[Lookup.scala 11:37]
  wire  _T_433 = _T_417 | _T_432; // @[Lookup.scala 11:37]
  wire  _T_434 = _T_413 | _T_433; // @[Lookup.scala 11:37]
  wire  _T_435 = _T_409 | _T_434; // @[Lookup.scala 11:37]
  wire  _T_436 = _T_405 | _T_435; // @[Lookup.scala 11:37]
  wire  _T_437 = _T_401 | _T_436; // @[Lookup.scala 11:37]
  wire  _T_438 = _T_397 | _T_437; // @[Lookup.scala 11:37]
  wire  _T_439 = _T_393 | _T_438; // @[Lookup.scala 11:37]
  wire  _T_440 = _T_389 | _T_439; // @[Lookup.scala 11:37]
  wire  _T_441 = _T_385 | _T_440; // @[Lookup.scala 11:37]
  wire  _T_442 = _T_381 | _T_441; // @[Lookup.scala 11:37]
  wire  _T_443 = _T_377 | _T_442; // @[Lookup.scala 11:37]
  wire  _T_444 = _T_373 | _T_443; // @[Lookup.scala 11:37]
  wire  _T_445 = _T_369 | _T_444; // @[Lookup.scala 11:37]
  wire  _T_446 = _T_365 | _T_445; // @[Lookup.scala 11:37]
  wire  _T_447 = _T_361 | _T_446; // @[Lookup.scala 11:37]
  wire  _T_448 = _T_357 | _T_447; // @[Lookup.scala 11:37]
  wire  _T_449 = _T_353 | _T_448; // @[Lookup.scala 11:37]
  wire  _T_450 = _T_349 | _T_449; // @[Lookup.scala 11:37]
  wire  _T_451 = _T_345 | _T_450; // @[Lookup.scala 11:37]
  wire  _T_452 = _T_341 | _T_451; // @[Lookup.scala 11:37]
  wire  _T_453 = _T_337 | _T_452; // @[Lookup.scala 11:37]
  wire  _T_454 = _T_333 | _T_453; // @[Lookup.scala 11:37]
  wire  _T_455 = _T_329 | _T_454; // @[Lookup.scala 11:37]
  wire  _T_456 = _T_325 | _T_455; // @[Lookup.scala 11:37]
  wire  _T_457 = _T_321 | _T_456; // @[Lookup.scala 11:37]
  wire  _T_458 = _T_317 | _T_457; // @[Lookup.scala 11:37]
  wire  _T_459 = _T_313 | _T_458; // @[Lookup.scala 11:37]
  wire  _T_460 = _T_309 | _T_459; // @[Lookup.scala 11:37]
  wire  _T_461 = _T_305 | _T_460; // @[Lookup.scala 11:37]
  wire  _T_462 = _T_301 | _T_461; // @[Lookup.scala 11:37]
  wire  _T_463 = _T_297 | _T_462; // @[Lookup.scala 11:37]
  wire  _T_464 = _T_293 | _T_463; // @[Lookup.scala 11:37]
  wire  _T_465 = _T_289 | _T_464; // @[Lookup.scala 11:37]
  wire  _T_466 = _T_285 | _T_465; // @[Lookup.scala 11:37]
  wire  _T_467 = _T_281 | _T_466; // @[Lookup.scala 11:37]
  wire  _T_468 = _T_277 | _T_467; // @[Lookup.scala 11:37]
  wire  _T_469 = _T_273 | _T_468; // @[Lookup.scala 11:37]
  wire  _T_470 = _T_269 | _T_469; // @[Lookup.scala 11:37]
  wire  _T_471 = _T_265 | _T_470; // @[Lookup.scala 11:37]
  wire  _T_472 = _T_261 | _T_471; // @[Lookup.scala 11:37]
  wire  _T_473 = _T_257 | _T_472; // @[Lookup.scala 11:37]
  wire  _T_474 = _T_253 | _T_473; // @[Lookup.scala 11:37]
  wire  _T_475 = _T_249 | _T_474; // @[Lookup.scala 11:37]
  wire  _T_476 = _T_245 | _T_475; // @[Lookup.scala 11:37]
  wire  _T_477 = _T_241 | _T_476; // @[Lookup.scala 11:37]
  wire  _T_478 = _T_237 | _T_477; // @[Lookup.scala 11:37]
  wire  cs_val_inst = _T_233 | _T_478; // @[Lookup.scala 11:37]
  wire [3:0] _T_492 = _T_377 ? 4'h6 : 4'h0; // @[Lookup.scala 11:37]
  wire [3:0] _T_493 = _T_373 ? 4'h5 : _T_492; // @[Lookup.scala 11:37]
  wire [3:0] _T_494 = _T_369 ? 4'h4 : _T_493; // @[Lookup.scala 11:37]
  wire [3:0] _T_495 = _T_365 ? 4'h3 : _T_494; // @[Lookup.scala 11:37]
  wire [3:0] _T_496 = _T_361 ? 4'h1 : _T_495; // @[Lookup.scala 11:37]
  wire [3:0] _T_497 = _T_357 ? 4'h2 : _T_496; // @[Lookup.scala 11:37]
  wire [3:0] _T_498 = _T_353 ? 4'h8 : _T_497; // @[Lookup.scala 11:37]
  wire [3:0] _T_499 = _T_349 ? 4'h7 : _T_498; // @[Lookup.scala 11:37]
  wire [3:0] _T_500 = _T_345 ? 4'h0 : _T_499; // @[Lookup.scala 11:37]
  wire [3:0] _T_501 = _T_341 ? 4'h0 : _T_500; // @[Lookup.scala 11:37]
  wire [3:0] _T_502 = _T_337 ? 4'h0 : _T_501; // @[Lookup.scala 11:37]
  wire [3:0] _T_503 = _T_333 ? 4'h0 : _T_502; // @[Lookup.scala 11:37]
  wire [3:0] _T_504 = _T_329 ? 4'h0 : _T_503; // @[Lookup.scala 11:37]
  wire [3:0] _T_505 = _T_325 ? 4'h0 : _T_504; // @[Lookup.scala 11:37]
  wire [3:0] _T_506 = _T_321 ? 4'h0 : _T_505; // @[Lookup.scala 11:37]
  wire [3:0] _T_507 = _T_317 ? 4'h0 : _T_506; // @[Lookup.scala 11:37]
  wire [3:0] _T_508 = _T_313 ? 4'h0 : _T_507; // @[Lookup.scala 11:37]
  wire [3:0] _T_509 = _T_309 ? 4'h0 : _T_508; // @[Lookup.scala 11:37]
  wire [3:0] _T_510 = _T_305 ? 4'h0 : _T_509; // @[Lookup.scala 11:37]
  wire [3:0] _T_511 = _T_301 ? 4'h0 : _T_510; // @[Lookup.scala 11:37]
  wire [3:0] _T_512 = _T_297 ? 4'h0 : _T_511; // @[Lookup.scala 11:37]
  wire [3:0] _T_513 = _T_293 ? 4'h0 : _T_512; // @[Lookup.scala 11:37]
  wire [3:0] _T_514 = _T_289 ? 4'h0 : _T_513; // @[Lookup.scala 11:37]
  wire [3:0] _T_515 = _T_285 ? 4'h0 : _T_514; // @[Lookup.scala 11:37]
  wire [3:0] _T_516 = _T_281 ? 4'h0 : _T_515; // @[Lookup.scala 11:37]
  wire [3:0] _T_517 = _T_277 ? 4'h0 : _T_516; // @[Lookup.scala 11:37]
  wire [3:0] _T_518 = _T_273 ? 4'h0 : _T_517; // @[Lookup.scala 11:37]
  wire [3:0] _T_519 = _T_269 ? 4'h0 : _T_518; // @[Lookup.scala 11:37]
  wire [3:0] _T_520 = _T_265 ? 4'h0 : _T_519; // @[Lookup.scala 11:37]
  wire [3:0] _T_521 = _T_261 ? 4'h0 : _T_520; // @[Lookup.scala 11:37]
  wire [3:0] _T_522 = _T_257 ? 4'h0 : _T_521; // @[Lookup.scala 11:37]
  wire [3:0] _T_523 = _T_253 ? 4'h0 : _T_522; // @[Lookup.scala 11:37]
  wire [3:0] _T_524 = _T_249 ? 4'h0 : _T_523; // @[Lookup.scala 11:37]
  wire [3:0] _T_525 = _T_245 ? 4'h0 : _T_524; // @[Lookup.scala 11:37]
  wire [3:0] _T_526 = _T_241 ? 4'h0 : _T_525; // @[Lookup.scala 11:37]
  wire [3:0] _T_527 = _T_237 ? 4'h0 : _T_526; // @[Lookup.scala 11:37]
  wire [1:0] _T_535 = _T_401 ? 2'h2 : 2'h0; // @[Lookup.scala 11:37]
  wire [1:0] _T_536 = _T_397 ? 2'h0 : _T_535; // @[Lookup.scala 11:37]
  wire [1:0] _T_537 = _T_393 ? 2'h0 : _T_536; // @[Lookup.scala 11:37]
  wire [1:0] _T_538 = _T_389 ? 2'h0 : _T_537; // @[Lookup.scala 11:37]
  wire [1:0] _T_539 = _T_385 ? 2'h2 : _T_538; // @[Lookup.scala 11:37]
  wire [1:0] _T_540 = _T_381 ? 2'h2 : _T_539; // @[Lookup.scala 11:37]
  wire [1:0] _T_541 = _T_377 ? 2'h0 : _T_540; // @[Lookup.scala 11:37]
  wire [1:0] _T_542 = _T_373 ? 2'h0 : _T_541; // @[Lookup.scala 11:37]
  wire [1:0] _T_543 = _T_369 ? 2'h0 : _T_542; // @[Lookup.scala 11:37]
  wire [1:0] _T_544 = _T_365 ? 2'h0 : _T_543; // @[Lookup.scala 11:37]
  wire [1:0] _T_545 = _T_361 ? 2'h0 : _T_544; // @[Lookup.scala 11:37]
  wire [1:0] _T_546 = _T_357 ? 2'h0 : _T_545; // @[Lookup.scala 11:37]
  wire [1:0] _T_547 = _T_353 ? 2'h0 : _T_546; // @[Lookup.scala 11:37]
  wire [1:0] _T_548 = _T_349 ? 2'h0 : _T_547; // @[Lookup.scala 11:37]
  wire [1:0] _T_549 = _T_345 ? 2'h0 : _T_548; // @[Lookup.scala 11:37]
  wire [1:0] _T_550 = _T_341 ? 2'h0 : _T_549; // @[Lookup.scala 11:37]
  wire [1:0] _T_551 = _T_337 ? 2'h0 : _T_550; // @[Lookup.scala 11:37]
  wire [1:0] _T_552 = _T_333 ? 2'h0 : _T_551; // @[Lookup.scala 11:37]
  wire [1:0] _T_553 = _T_329 ? 2'h0 : _T_552; // @[Lookup.scala 11:37]
  wire [1:0] _T_554 = _T_325 ? 2'h0 : _T_553; // @[Lookup.scala 11:37]
  wire [1:0] _T_555 = _T_321 ? 2'h0 : _T_554; // @[Lookup.scala 11:37]
  wire [1:0] _T_556 = _T_317 ? 2'h0 : _T_555; // @[Lookup.scala 11:37]
  wire [1:0] _T_557 = _T_313 ? 2'h0 : _T_556; // @[Lookup.scala 11:37]
  wire [1:0] _T_558 = _T_309 ? 2'h0 : _T_557; // @[Lookup.scala 11:37]
  wire [1:0] _T_559 = _T_305 ? 2'h0 : _T_558; // @[Lookup.scala 11:37]
  wire [1:0] _T_560 = _T_301 ? 2'h0 : _T_559; // @[Lookup.scala 11:37]
  wire [1:0] _T_561 = _T_297 ? 2'h0 : _T_560; // @[Lookup.scala 11:37]
  wire [1:0] _T_562 = _T_293 ? 2'h0 : _T_561; // @[Lookup.scala 11:37]
  wire [1:0] _T_563 = _T_289 ? 2'h0 : _T_562; // @[Lookup.scala 11:37]
  wire [1:0] _T_564 = _T_285 ? 2'h0 : _T_563; // @[Lookup.scala 11:37]
  wire [1:0] _T_565 = _T_281 ? 2'h0 : _T_564; // @[Lookup.scala 11:37]
  wire [1:0] _T_566 = _T_277 ? 2'h0 : _T_565; // @[Lookup.scala 11:37]
  wire [1:0] _T_567 = _T_273 ? 2'h0 : _T_566; // @[Lookup.scala 11:37]
  wire [1:0] _T_568 = _T_269 ? 2'h0 : _T_567; // @[Lookup.scala 11:37]
  wire [1:0] _T_569 = _T_265 ? 2'h1 : _T_568; // @[Lookup.scala 11:37]
  wire [1:0] _T_570 = _T_261 ? 2'h0 : _T_569; // @[Lookup.scala 11:37]
  wire [1:0] _T_571 = _T_257 ? 2'h0 : _T_570; // @[Lookup.scala 11:37]
  wire [1:0] _T_572 = _T_253 ? 2'h0 : _T_571; // @[Lookup.scala 11:37]
  wire [1:0] _T_573 = _T_249 ? 2'h0 : _T_572; // @[Lookup.scala 11:37]
  wire [1:0] _T_574 = _T_245 ? 2'h0 : _T_573; // @[Lookup.scala 11:37]
  wire [1:0] _T_575 = _T_241 ? 2'h0 : _T_574; // @[Lookup.scala 11:37]
  wire [1:0] _T_576 = _T_237 ? 2'h0 : _T_575; // @[Lookup.scala 11:37]
  wire [2:0] _T_590 = _T_377 ? 3'h3 : 3'h0; // @[Lookup.scala 11:37]
  wire [2:0] _T_591 = _T_373 ? 3'h3 : _T_590; // @[Lookup.scala 11:37]
  wire [2:0] _T_592 = _T_369 ? 3'h3 : _T_591; // @[Lookup.scala 11:37]
  wire [2:0] _T_593 = _T_365 ? 3'h3 : _T_592; // @[Lookup.scala 11:37]
  wire [2:0] _T_594 = _T_361 ? 3'h3 : _T_593; // @[Lookup.scala 11:37]
  wire [2:0] _T_595 = _T_357 ? 3'h3 : _T_594; // @[Lookup.scala 11:37]
  wire [2:0] _T_596 = _T_353 ? 3'h1 : _T_595; // @[Lookup.scala 11:37]
  wire [2:0] _T_597 = _T_349 ? 3'h5 : _T_596; // @[Lookup.scala 11:37]
  wire [2:0] _T_598 = _T_345 ? 3'h0 : _T_597; // @[Lookup.scala 11:37]
  wire [2:0] _T_599 = _T_341 ? 3'h0 : _T_598; // @[Lookup.scala 11:37]
  wire [2:0] _T_600 = _T_337 ? 3'h0 : _T_599; // @[Lookup.scala 11:37]
  wire [2:0] _T_601 = _T_333 ? 3'h0 : _T_600; // @[Lookup.scala 11:37]
  wire [2:0] _T_602 = _T_329 ? 3'h0 : _T_601; // @[Lookup.scala 11:37]
  wire [2:0] _T_603 = _T_325 ? 3'h0 : _T_602; // @[Lookup.scala 11:37]
  wire [2:0] _T_604 = _T_321 ? 3'h0 : _T_603; // @[Lookup.scala 11:37]
  wire [2:0] _T_605 = _T_317 ? 3'h0 : _T_604; // @[Lookup.scala 11:37]
  wire [2:0] _T_606 = _T_313 ? 3'h0 : _T_605; // @[Lookup.scala 11:37]
  wire [2:0] _T_607 = _T_309 ? 3'h0 : _T_606; // @[Lookup.scala 11:37]
  wire [2:0] _T_608 = _T_305 ? 3'h1 : _T_607; // @[Lookup.scala 11:37]
  wire [2:0] _T_609 = _T_301 ? 3'h1 : _T_608; // @[Lookup.scala 11:37]
  wire [2:0] _T_610 = _T_297 ? 3'h1 : _T_609; // @[Lookup.scala 11:37]
  wire [2:0] _T_611 = _T_293 ? 3'h1 : _T_610; // @[Lookup.scala 11:37]
  wire [2:0] _T_612 = _T_289 ? 3'h1 : _T_611; // @[Lookup.scala 11:37]
  wire [2:0] _T_613 = _T_285 ? 3'h1 : _T_612; // @[Lookup.scala 11:37]
  wire [2:0] _T_614 = _T_281 ? 3'h1 : _T_613; // @[Lookup.scala 11:37]
  wire [2:0] _T_615 = _T_277 ? 3'h1 : _T_614; // @[Lookup.scala 11:37]
  wire [2:0] _T_616 = _T_273 ? 3'h1 : _T_615; // @[Lookup.scala 11:37]
  wire [2:0] _T_617 = _T_269 ? 3'h4 : _T_616; // @[Lookup.scala 11:37]
  wire [2:0] _T_618 = _T_265 ? 3'h4 : _T_617; // @[Lookup.scala 11:37]
  wire [2:0] _T_619 = _T_261 ? 3'h2 : _T_618; // @[Lookup.scala 11:37]
  wire [2:0] _T_620 = _T_257 ? 3'h2 : _T_619; // @[Lookup.scala 11:37]
  wire [2:0] _T_621 = _T_253 ? 3'h2 : _T_620; // @[Lookup.scala 11:37]
  wire [2:0] _T_622 = _T_249 ? 3'h1 : _T_621; // @[Lookup.scala 11:37]
  wire [2:0] _T_623 = _T_245 ? 3'h1 : _T_622; // @[Lookup.scala 11:37]
  wire [2:0] _T_624 = _T_241 ? 3'h1 : _T_623; // @[Lookup.scala 11:37]
  wire [2:0] _T_625 = _T_237 ? 3'h1 : _T_624; // @[Lookup.scala 11:37]
  wire  _T_634 = _T_397 | _T_401; // @[Lookup.scala 11:37]
  wire  _T_635 = _T_393 | _T_634; // @[Lookup.scala 11:37]
  wire  _T_636 = _T_389 | _T_635; // @[Lookup.scala 11:37]
  wire  _T_637 = _T_385 | _T_636; // @[Lookup.scala 11:37]
  wire  _T_638 = _T_381 | _T_637; // @[Lookup.scala 11:37]
  wire  _T_639 = _T_377 | _T_638; // @[Lookup.scala 11:37]
  wire  _T_640 = _T_373 | _T_639; // @[Lookup.scala 11:37]
  wire  _T_641 = _T_369 | _T_640; // @[Lookup.scala 11:37]
  wire  _T_642 = _T_365 | _T_641; // @[Lookup.scala 11:37]
  wire  _T_643 = _T_361 | _T_642; // @[Lookup.scala 11:37]
  wire  _T_644 = _T_357 | _T_643; // @[Lookup.scala 11:37]
  wire  _T_645 = _T_353 | _T_644; // @[Lookup.scala 11:37]
  wire  _T_646 = _T_349 ? 1'h0 : _T_645; // @[Lookup.scala 11:37]
  wire  _T_647 = _T_345 | _T_646; // @[Lookup.scala 11:37]
  wire  _T_648 = _T_341 | _T_647; // @[Lookup.scala 11:37]
  wire  _T_649 = _T_337 | _T_648; // @[Lookup.scala 11:37]
  wire  _T_650 = _T_333 | _T_649; // @[Lookup.scala 11:37]
  wire  _T_651 = _T_329 | _T_650; // @[Lookup.scala 11:37]
  wire  _T_652 = _T_325 | _T_651; // @[Lookup.scala 11:37]
  wire  _T_653 = _T_321 | _T_652; // @[Lookup.scala 11:37]
  wire  _T_654 = _T_317 | _T_653; // @[Lookup.scala 11:37]
  wire  _T_655 = _T_313 | _T_654; // @[Lookup.scala 11:37]
  wire  _T_656 = _T_309 | _T_655; // @[Lookup.scala 11:37]
  wire  _T_657 = _T_305 | _T_656; // @[Lookup.scala 11:37]
  wire  _T_658 = _T_301 | _T_657; // @[Lookup.scala 11:37]
  wire  _T_659 = _T_297 | _T_658; // @[Lookup.scala 11:37]
  wire  _T_660 = _T_293 | _T_659; // @[Lookup.scala 11:37]
  wire  _T_661 = _T_289 | _T_660; // @[Lookup.scala 11:37]
  wire  _T_662 = _T_285 | _T_661; // @[Lookup.scala 11:37]
  wire  _T_663 = _T_281 | _T_662; // @[Lookup.scala 11:37]
  wire  _T_664 = _T_277 | _T_663; // @[Lookup.scala 11:37]
  wire  _T_665 = _T_273 | _T_664; // @[Lookup.scala 11:37]
  wire  _T_666 = _T_269 ? 1'h0 : _T_665; // @[Lookup.scala 11:37]
  wire  _T_667 = _T_265 ? 1'h0 : _T_666; // @[Lookup.scala 11:37]
  wire  _T_668 = _T_261 | _T_667; // @[Lookup.scala 11:37]
  wire  _T_669 = _T_257 | _T_668; // @[Lookup.scala 11:37]
  wire  _T_670 = _T_253 | _T_669; // @[Lookup.scala 11:37]
  wire  _T_671 = _T_249 | _T_670; // @[Lookup.scala 11:37]
  wire  _T_672 = _T_245 | _T_671; // @[Lookup.scala 11:37]
  wire  _T_673 = _T_241 | _T_672; // @[Lookup.scala 11:37]
  wire  _T_674 = _T_237 | _T_673; // @[Lookup.scala 11:37]
  wire  cs_rs1_oen = _T_233 | _T_674; // @[Lookup.scala 11:37]
  wire  _T_694 = _T_353 ? 1'h0 : _T_644; // @[Lookup.scala 11:37]
  wire  _T_695 = _T_349 ? 1'h0 : _T_694; // @[Lookup.scala 11:37]
  wire  _T_696 = _T_345 | _T_695; // @[Lookup.scala 11:37]
  wire  _T_697 = _T_341 | _T_696; // @[Lookup.scala 11:37]
  wire  _T_698 = _T_337 | _T_697; // @[Lookup.scala 11:37]
  wire  _T_699 = _T_333 | _T_698; // @[Lookup.scala 11:37]
  wire  _T_700 = _T_329 | _T_699; // @[Lookup.scala 11:37]
  wire  _T_701 = _T_325 | _T_700; // @[Lookup.scala 11:37]
  wire  _T_702 = _T_321 | _T_701; // @[Lookup.scala 11:37]
  wire  _T_703 = _T_317 | _T_702; // @[Lookup.scala 11:37]
  wire  _T_704 = _T_313 | _T_703; // @[Lookup.scala 11:37]
  wire  _T_705 = _T_309 | _T_704; // @[Lookup.scala 11:37]
  wire  _T_706 = _T_305 ? 1'h0 : _T_705; // @[Lookup.scala 11:37]
  wire  _T_707 = _T_301 ? 1'h0 : _T_706; // @[Lookup.scala 11:37]
  wire  _T_708 = _T_297 ? 1'h0 : _T_707; // @[Lookup.scala 11:37]
  wire  _T_709 = _T_293 ? 1'h0 : _T_708; // @[Lookup.scala 11:37]
  wire  _T_710 = _T_289 ? 1'h0 : _T_709; // @[Lookup.scala 11:37]
  wire  _T_711 = _T_285 ? 1'h0 : _T_710; // @[Lookup.scala 11:37]
  wire  _T_712 = _T_281 ? 1'h0 : _T_711; // @[Lookup.scala 11:37]
  wire  _T_713 = _T_277 ? 1'h0 : _T_712; // @[Lookup.scala 11:37]
  wire  _T_714 = _T_273 ? 1'h0 : _T_713; // @[Lookup.scala 11:37]
  wire  _T_715 = _T_269 ? 1'h0 : _T_714; // @[Lookup.scala 11:37]
  wire  _T_716 = _T_265 ? 1'h0 : _T_715; // @[Lookup.scala 11:37]
  wire  _T_717 = _T_261 | _T_716; // @[Lookup.scala 11:37]
  wire  _T_718 = _T_257 | _T_717; // @[Lookup.scala 11:37]
  wire  _T_719 = _T_253 | _T_718; // @[Lookup.scala 11:37]
  wire  _T_720 = _T_249 ? 1'h0 : _T_719; // @[Lookup.scala 11:37]
  wire  _T_721 = _T_245 ? 1'h0 : _T_720; // @[Lookup.scala 11:37]
  wire  _T_722 = _T_241 ? 1'h0 : _T_721; // @[Lookup.scala 11:37]
  wire  _T_723 = _T_237 ? 1'h0 : _T_722; // @[Lookup.scala 11:37]
  wire  cs_rs2_oen = _T_233 ? 1'h0 : _T_723; // @[Lookup.scala 11:37]
  wire [3:0] _T_731 = _T_401 ? 4'ha : 4'h0; // @[Lookup.scala 11:37]
  wire [3:0] _T_732 = _T_397 ? 4'ha : _T_731; // @[Lookup.scala 11:37]
  wire [3:0] _T_733 = _T_393 ? 4'ha : _T_732; // @[Lookup.scala 11:37]
  wire [3:0] _T_734 = _T_389 ? 4'ha : _T_733; // @[Lookup.scala 11:37]
  wire [3:0] _T_735 = _T_385 ? 4'ha : _T_734; // @[Lookup.scala 11:37]
  wire [3:0] _T_736 = _T_381 ? 4'ha : _T_735; // @[Lookup.scala 11:37]
  wire [3:0] _T_737 = _T_377 ? 4'h0 : _T_736; // @[Lookup.scala 11:37]
  wire [3:0] _T_738 = _T_373 ? 4'h0 : _T_737; // @[Lookup.scala 11:37]
  wire [3:0] _T_739 = _T_369 ? 4'h0 : _T_738; // @[Lookup.scala 11:37]
  wire [3:0] _T_740 = _T_365 ? 4'h0 : _T_739; // @[Lookup.scala 11:37]
  wire [3:0] _T_741 = _T_361 ? 4'h0 : _T_740; // @[Lookup.scala 11:37]
  wire [3:0] _T_742 = _T_357 ? 4'h0 : _T_741; // @[Lookup.scala 11:37]
  wire [3:0] _T_743 = _T_353 ? 4'h0 : _T_742; // @[Lookup.scala 11:37]
  wire [3:0] _T_744 = _T_349 ? 4'h0 : _T_743; // @[Lookup.scala 11:37]
  wire [3:0] _T_745 = _T_345 ? 4'h3 : _T_744; // @[Lookup.scala 11:37]
  wire [3:0] _T_746 = _T_341 ? 4'h4 : _T_745; // @[Lookup.scala 11:37]
  wire [3:0] _T_747 = _T_337 ? 4'h7 : _T_746; // @[Lookup.scala 11:37]
  wire [3:0] _T_748 = _T_333 ? 4'h6 : _T_747; // @[Lookup.scala 11:37]
  wire [3:0] _T_749 = _T_329 ? 4'h5 : _T_748; // @[Lookup.scala 11:37]
  wire [3:0] _T_750 = _T_325 ? 4'h9 : _T_749; // @[Lookup.scala 11:37]
  wire [3:0] _T_751 = _T_321 ? 4'h8 : _T_750; // @[Lookup.scala 11:37]
  wire [3:0] _T_752 = _T_317 ? 4'h1 : _T_751; // @[Lookup.scala 11:37]
  wire [3:0] _T_753 = _T_313 ? 4'h0 : _T_752; // @[Lookup.scala 11:37]
  wire [3:0] _T_754 = _T_309 ? 4'h2 : _T_753; // @[Lookup.scala 11:37]
  wire [3:0] _T_755 = _T_305 ? 4'h3 : _T_754; // @[Lookup.scala 11:37]
  wire [3:0] _T_756 = _T_301 ? 4'h4 : _T_755; // @[Lookup.scala 11:37]
  wire [3:0] _T_757 = _T_297 ? 4'h2 : _T_756; // @[Lookup.scala 11:37]
  wire [3:0] _T_758 = _T_293 ? 4'h9 : _T_757; // @[Lookup.scala 11:37]
  wire [3:0] _T_759 = _T_289 ? 4'h8 : _T_758; // @[Lookup.scala 11:37]
  wire [3:0] _T_760 = _T_285 ? 4'h7 : _T_759; // @[Lookup.scala 11:37]
  wire [3:0] _T_761 = _T_281 ? 4'h6 : _T_760; // @[Lookup.scala 11:37]
  wire [3:0] _T_762 = _T_277 ? 4'h5 : _T_761; // @[Lookup.scala 11:37]
  wire [3:0] _T_763 = _T_273 ? 4'h0 : _T_762; // @[Lookup.scala 11:37]
  wire [3:0] _T_764 = _T_269 ? 4'hb : _T_763; // @[Lookup.scala 11:37]
  wire [3:0] _T_765 = _T_265 ? 4'h0 : _T_764; // @[Lookup.scala 11:37]
  wire [3:0] _T_766 = _T_261 ? 4'h0 : _T_765; // @[Lookup.scala 11:37]
  wire [3:0] _T_767 = _T_257 ? 4'h0 : _T_766; // @[Lookup.scala 11:37]
  wire [3:0] _T_768 = _T_253 ? 4'h0 : _T_767; // @[Lookup.scala 11:37]
  wire [3:0] _T_769 = _T_249 ? 4'h0 : _T_768; // @[Lookup.scala 11:37]
  wire [3:0] _T_770 = _T_245 ? 4'h0 : _T_769; // @[Lookup.scala 11:37]
  wire [3:0] _T_771 = _T_241 ? 4'h0 : _T_770; // @[Lookup.scala 11:37]
  wire [3:0] _T_772 = _T_237 ? 4'h0 : _T_771; // @[Lookup.scala 11:37]
  wire [1:0] _T_780 = _T_401 ? 2'h3 : 2'h0; // @[Lookup.scala 11:37]
  wire [1:0] _T_781 = _T_397 ? 2'h3 : _T_780; // @[Lookup.scala 11:37]
  wire [1:0] _T_782 = _T_393 ? 2'h3 : _T_781; // @[Lookup.scala 11:37]
  wire [1:0] _T_783 = _T_389 ? 2'h3 : _T_782; // @[Lookup.scala 11:37]
  wire [1:0] _T_784 = _T_385 ? 2'h3 : _T_783; // @[Lookup.scala 11:37]
  wire [1:0] _T_785 = _T_381 ? 2'h3 : _T_784; // @[Lookup.scala 11:37]
  wire [1:0] _T_786 = _T_377 ? 2'h0 : _T_785; // @[Lookup.scala 11:37]
  wire [1:0] _T_787 = _T_373 ? 2'h0 : _T_786; // @[Lookup.scala 11:37]
  wire [1:0] _T_788 = _T_369 ? 2'h0 : _T_787; // @[Lookup.scala 11:37]
  wire [1:0] _T_789 = _T_365 ? 2'h0 : _T_788; // @[Lookup.scala 11:37]
  wire [1:0] _T_790 = _T_361 ? 2'h0 : _T_789; // @[Lookup.scala 11:37]
  wire [1:0] _T_791 = _T_357 ? 2'h0 : _T_790; // @[Lookup.scala 11:37]
  wire [1:0] _T_792 = _T_353 ? 2'h2 : _T_791; // @[Lookup.scala 11:37]
  wire [1:0] _T_793 = _T_349 ? 2'h2 : _T_792; // @[Lookup.scala 11:37]
  wire [1:0] _T_794 = _T_345 ? 2'h0 : _T_793; // @[Lookup.scala 11:37]
  wire [1:0] _T_795 = _T_341 ? 2'h0 : _T_794; // @[Lookup.scala 11:37]
  wire [1:0] _T_796 = _T_337 ? 2'h0 : _T_795; // @[Lookup.scala 11:37]
  wire [1:0] _T_797 = _T_333 ? 2'h0 : _T_796; // @[Lookup.scala 11:37]
  wire [1:0] _T_798 = _T_329 ? 2'h0 : _T_797; // @[Lookup.scala 11:37]
  wire [1:0] _T_799 = _T_325 ? 2'h0 : _T_798; // @[Lookup.scala 11:37]
  wire [1:0] _T_800 = _T_321 ? 2'h0 : _T_799; // @[Lookup.scala 11:37]
  wire [1:0] _T_801 = _T_317 ? 2'h0 : _T_800; // @[Lookup.scala 11:37]
  wire [1:0] _T_802 = _T_313 ? 2'h0 : _T_801; // @[Lookup.scala 11:37]
  wire [1:0] _T_803 = _T_309 ? 2'h0 : _T_802; // @[Lookup.scala 11:37]
  wire [1:0] _T_804 = _T_305 ? 2'h0 : _T_803; // @[Lookup.scala 11:37]
  wire [1:0] _T_805 = _T_301 ? 2'h0 : _T_804; // @[Lookup.scala 11:37]
  wire [1:0] _T_806 = _T_297 ? 2'h0 : _T_805; // @[Lookup.scala 11:37]
  wire [1:0] _T_807 = _T_293 ? 2'h0 : _T_806; // @[Lookup.scala 11:37]
  wire [1:0] _T_808 = _T_289 ? 2'h0 : _T_807; // @[Lookup.scala 11:37]
  wire [1:0] _T_809 = _T_285 ? 2'h0 : _T_808; // @[Lookup.scala 11:37]
  wire [1:0] _T_810 = _T_281 ? 2'h0 : _T_809; // @[Lookup.scala 11:37]
  wire [1:0] _T_811 = _T_277 ? 2'h0 : _T_810; // @[Lookup.scala 11:37]
  wire [1:0] _T_812 = _T_273 ? 2'h0 : _T_811; // @[Lookup.scala 11:37]
  wire [1:0] _T_813 = _T_269 ? 2'h0 : _T_812; // @[Lookup.scala 11:37]
  wire [1:0] _T_814 = _T_265 ? 2'h0 : _T_813; // @[Lookup.scala 11:37]
  wire [1:0] _T_815 = _T_261 ? 2'h0 : _T_814; // @[Lookup.scala 11:37]
  wire [1:0] _T_816 = _T_257 ? 2'h0 : _T_815; // @[Lookup.scala 11:37]
  wire [1:0] _T_817 = _T_253 ? 2'h0 : _T_816; // @[Lookup.scala 11:37]
  wire [1:0] _T_818 = _T_249 ? 2'h1 : _T_817; // @[Lookup.scala 11:37]
  wire [1:0] _T_819 = _T_245 ? 2'h1 : _T_818; // @[Lookup.scala 11:37]
  wire [1:0] _T_820 = _T_241 ? 2'h1 : _T_819; // @[Lookup.scala 11:37]
  wire [1:0] _T_821 = _T_237 ? 2'h1 : _T_820; // @[Lookup.scala 11:37]
  wire  _T_835 = _T_377 ? 1'h0 : _T_638; // @[Lookup.scala 11:37]
  wire  _T_836 = _T_373 ? 1'h0 : _T_835; // @[Lookup.scala 11:37]
  wire  _T_837 = _T_369 ? 1'h0 : _T_836; // @[Lookup.scala 11:37]
  wire  _T_838 = _T_365 ? 1'h0 : _T_837; // @[Lookup.scala 11:37]
  wire  _T_839 = _T_361 ? 1'h0 : _T_838; // @[Lookup.scala 11:37]
  wire  _T_840 = _T_357 ? 1'h0 : _T_839; // @[Lookup.scala 11:37]
  wire  _T_841 = _T_353 | _T_840; // @[Lookup.scala 11:37]
  wire  _T_842 = _T_349 | _T_841; // @[Lookup.scala 11:37]
  wire  _T_843 = _T_345 | _T_842; // @[Lookup.scala 11:37]
  wire  _T_844 = _T_341 | _T_843; // @[Lookup.scala 11:37]
  wire  _T_845 = _T_337 | _T_844; // @[Lookup.scala 11:37]
  wire  _T_846 = _T_333 | _T_845; // @[Lookup.scala 11:37]
  wire  _T_847 = _T_329 | _T_846; // @[Lookup.scala 11:37]
  wire  _T_848 = _T_325 | _T_847; // @[Lookup.scala 11:37]
  wire  _T_849 = _T_321 | _T_848; // @[Lookup.scala 11:37]
  wire  _T_850 = _T_317 | _T_849; // @[Lookup.scala 11:37]
  wire  _T_851 = _T_313 | _T_850; // @[Lookup.scala 11:37]
  wire  _T_852 = _T_309 | _T_851; // @[Lookup.scala 11:37]
  wire  _T_853 = _T_305 | _T_852; // @[Lookup.scala 11:37]
  wire  _T_854 = _T_301 | _T_853; // @[Lookup.scala 11:37]
  wire  _T_855 = _T_297 | _T_854; // @[Lookup.scala 11:37]
  wire  _T_856 = _T_293 | _T_855; // @[Lookup.scala 11:37]
  wire  _T_857 = _T_289 | _T_856; // @[Lookup.scala 11:37]
  wire  _T_858 = _T_285 | _T_857; // @[Lookup.scala 11:37]
  wire  _T_859 = _T_281 | _T_858; // @[Lookup.scala 11:37]
  wire  _T_860 = _T_277 | _T_859; // @[Lookup.scala 11:37]
  wire  _T_861 = _T_273 | _T_860; // @[Lookup.scala 11:37]
  wire  _T_862 = _T_269 | _T_861; // @[Lookup.scala 11:37]
  wire  _T_863 = _T_265 | _T_862; // @[Lookup.scala 11:37]
  wire  _T_864 = _T_261 ? 1'h0 : _T_863; // @[Lookup.scala 11:37]
  wire  _T_865 = _T_257 ? 1'h0 : _T_864; // @[Lookup.scala 11:37]
  wire  _T_866 = _T_253 ? 1'h0 : _T_865; // @[Lookup.scala 11:37]
  wire  _T_867 = _T_249 | _T_866; // @[Lookup.scala 11:37]
  wire  _T_868 = _T_245 | _T_867; // @[Lookup.scala 11:37]
  wire  _T_869 = _T_241 | _T_868; // @[Lookup.scala 11:37]
  wire  _T_870 = _T_237 | _T_869; // @[Lookup.scala 11:37]
  wire  _T_872 = _T_425 ? 1'h0 : _T_429; // @[Lookup.scala 11:37]
  wire  _T_873 = _T_421 ? 1'h0 : _T_872; // @[Lookup.scala 11:37]
  wire  _T_874 = _T_417 ? 1'h0 : _T_873; // @[Lookup.scala 11:37]
  wire  _T_875 = _T_413 ? 1'h0 : _T_874; // @[Lookup.scala 11:37]
  wire  _T_876 = _T_409 ? 1'h0 : _T_875; // @[Lookup.scala 11:37]
  wire  _T_877 = _T_405 ? 1'h0 : _T_876; // @[Lookup.scala 11:37]
  wire  _T_878 = _T_401 ? 1'h0 : _T_877; // @[Lookup.scala 11:37]
  wire  _T_879 = _T_397 ? 1'h0 : _T_878; // @[Lookup.scala 11:37]
  wire  _T_880 = _T_393 ? 1'h0 : _T_879; // @[Lookup.scala 11:37]
  wire  _T_881 = _T_389 ? 1'h0 : _T_880; // @[Lookup.scala 11:37]
  wire  _T_882 = _T_385 ? 1'h0 : _T_881; // @[Lookup.scala 11:37]
  wire  _T_883 = _T_381 ? 1'h0 : _T_882; // @[Lookup.scala 11:37]
  wire  _T_884 = _T_377 ? 1'h0 : _T_883; // @[Lookup.scala 11:37]
  wire  _T_885 = _T_373 ? 1'h0 : _T_884; // @[Lookup.scala 11:37]
  wire  _T_886 = _T_369 ? 1'h0 : _T_885; // @[Lookup.scala 11:37]
  wire  _T_887 = _T_365 ? 1'h0 : _T_886; // @[Lookup.scala 11:37]
  wire  _T_888 = _T_361 ? 1'h0 : _T_887; // @[Lookup.scala 11:37]
  wire  _T_889 = _T_357 ? 1'h0 : _T_888; // @[Lookup.scala 11:37]
  wire  _T_890 = _T_353 ? 1'h0 : _T_889; // @[Lookup.scala 11:37]
  wire  _T_891 = _T_349 ? 1'h0 : _T_890; // @[Lookup.scala 11:37]
  wire  _T_892 = _T_345 ? 1'h0 : _T_891; // @[Lookup.scala 11:37]
  wire  _T_893 = _T_341 ? 1'h0 : _T_892; // @[Lookup.scala 11:37]
  wire  _T_894 = _T_337 ? 1'h0 : _T_893; // @[Lookup.scala 11:37]
  wire  _T_895 = _T_333 ? 1'h0 : _T_894; // @[Lookup.scala 11:37]
  wire  _T_896 = _T_329 ? 1'h0 : _T_895; // @[Lookup.scala 11:37]
  wire  _T_897 = _T_325 ? 1'h0 : _T_896; // @[Lookup.scala 11:37]
  wire  _T_898 = _T_321 ? 1'h0 : _T_897; // @[Lookup.scala 11:37]
  wire  _T_899 = _T_317 ? 1'h0 : _T_898; // @[Lookup.scala 11:37]
  wire  _T_900 = _T_313 ? 1'h0 : _T_899; // @[Lookup.scala 11:37]
  wire  _T_901 = _T_309 ? 1'h0 : _T_900; // @[Lookup.scala 11:37]
  wire  _T_902 = _T_305 ? 1'h0 : _T_901; // @[Lookup.scala 11:37]
  wire  _T_903 = _T_301 ? 1'h0 : _T_902; // @[Lookup.scala 11:37]
  wire  _T_904 = _T_297 ? 1'h0 : _T_903; // @[Lookup.scala 11:37]
  wire  _T_905 = _T_293 ? 1'h0 : _T_904; // @[Lookup.scala 11:37]
  wire  _T_906 = _T_289 ? 1'h0 : _T_905; // @[Lookup.scala 11:37]
  wire  _T_907 = _T_285 ? 1'h0 : _T_906; // @[Lookup.scala 11:37]
  wire  _T_908 = _T_281 ? 1'h0 : _T_907; // @[Lookup.scala 11:37]
  wire  _T_909 = _T_277 ? 1'h0 : _T_908; // @[Lookup.scala 11:37]
  wire  _T_910 = _T_273 ? 1'h0 : _T_909; // @[Lookup.scala 11:37]
  wire  _T_911 = _T_269 ? 1'h0 : _T_910; // @[Lookup.scala 11:37]
  wire  _T_912 = _T_265 ? 1'h0 : _T_911; // @[Lookup.scala 11:37]
  wire  _T_913 = _T_261 | _T_912; // @[Lookup.scala 11:37]
  wire  _T_914 = _T_257 | _T_913; // @[Lookup.scala 11:37]
  wire  _T_915 = _T_253 | _T_914; // @[Lookup.scala 11:37]
  wire  _T_916 = _T_249 | _T_915; // @[Lookup.scala 11:37]
  wire  _T_917 = _T_245 | _T_916; // @[Lookup.scala 11:37]
  wire  _T_918 = _T_241 | _T_917; // @[Lookup.scala 11:37]
  wire  _T_919 = _T_237 | _T_918; // @[Lookup.scala 11:37]
  wire  cs0_3 = _T_233 | _T_919; // @[Lookup.scala 11:37]
  wire  _T_963 = _T_257 | _T_261; // @[Lookup.scala 11:37]
  wire  _T_964 = _T_253 | _T_963; // @[Lookup.scala 11:37]
  wire  _T_965 = _T_249 ? 1'h0 : _T_964; // @[Lookup.scala 11:37]
  wire  _T_966 = _T_245 ? 1'h0 : _T_965; // @[Lookup.scala 11:37]
  wire  _T_967 = _T_241 ? 1'h0 : _T_966; // @[Lookup.scala 11:37]
  wire  _T_968 = _T_237 ? 1'h0 : _T_967; // @[Lookup.scala 11:37]
  wire  cs0_4 = _T_233 ? 1'h0 : _T_968; // @[Lookup.scala 11:37]
  wire [2:0] _T_1011 = _T_261 ? 3'h2 : 3'h0; // @[Lookup.scala 11:37]
  wire [2:0] _T_1012 = _T_257 ? 3'h1 : _T_1011; // @[Lookup.scala 11:37]
  wire [2:0] _T_1013 = _T_253 ? 3'h3 : _T_1012; // @[Lookup.scala 11:37]
  wire [2:0] _T_1014 = _T_249 ? 3'h6 : _T_1013; // @[Lookup.scala 11:37]
  wire [2:0] _T_1015 = _T_245 ? 3'h2 : _T_1014; // @[Lookup.scala 11:37]
  wire [2:0] _T_1016 = _T_241 ? 3'h5 : _T_1015; // @[Lookup.scala 11:37]
  wire [2:0] _T_1017 = _T_237 ? 3'h1 : _T_1016; // @[Lookup.scala 11:37]
  wire [2:0] _T_1021 = _T_417 ? 3'h4 : 3'h0; // @[Lookup.scala 11:37]
  wire [2:0] _T_1022 = _T_413 ? 3'h4 : _T_1021; // @[Lookup.scala 11:37]
  wire [2:0] _T_1023 = _T_409 ? 3'h4 : _T_1022; // @[Lookup.scala 11:37]
  wire [2:0] _T_1024 = _T_405 ? 3'h4 : _T_1023; // @[Lookup.scala 11:37]
  wire [2:0] _T_1025 = _T_401 ? 3'h3 : _T_1024; // @[Lookup.scala 11:37]
  wire [2:0] _T_1026 = _T_397 ? 3'h3 : _T_1025; // @[Lookup.scala 11:37]
  wire [2:0] _T_1027 = _T_393 ? 3'h2 : _T_1026; // @[Lookup.scala 11:37]
  wire [2:0] _T_1028 = _T_389 ? 3'h1 : _T_1027; // @[Lookup.scala 11:37]
  wire [2:0] _T_1029 = _T_385 ? 3'h2 : _T_1028; // @[Lookup.scala 11:37]
  wire [2:0] _T_1030 = _T_381 ? 3'h1 : _T_1029; // @[Lookup.scala 11:37]
  wire [2:0] _T_1031 = _T_377 ? 3'h0 : _T_1030; // @[Lookup.scala 11:37]
  wire [2:0] _T_1032 = _T_373 ? 3'h0 : _T_1031; // @[Lookup.scala 11:37]
  wire [2:0] _T_1033 = _T_369 ? 3'h0 : _T_1032; // @[Lookup.scala 11:37]
  wire [2:0] _T_1034 = _T_365 ? 3'h0 : _T_1033; // @[Lookup.scala 11:37]
  wire [2:0] _T_1035 = _T_361 ? 3'h0 : _T_1034; // @[Lookup.scala 11:37]
  wire [2:0] _T_1036 = _T_357 ? 3'h0 : _T_1035; // @[Lookup.scala 11:37]
  wire [2:0] _T_1037 = _T_353 ? 3'h0 : _T_1036; // @[Lookup.scala 11:37]
  wire [2:0] _T_1038 = _T_349 ? 3'h0 : _T_1037; // @[Lookup.scala 11:37]
  wire [2:0] _T_1039 = _T_345 ? 3'h0 : _T_1038; // @[Lookup.scala 11:37]
  wire [2:0] _T_1040 = _T_341 ? 3'h0 : _T_1039; // @[Lookup.scala 11:37]
  wire [2:0] _T_1041 = _T_337 ? 3'h0 : _T_1040; // @[Lookup.scala 11:37]
  wire [2:0] _T_1042 = _T_333 ? 3'h0 : _T_1041; // @[Lookup.scala 11:37]
  wire [2:0] _T_1043 = _T_329 ? 3'h0 : _T_1042; // @[Lookup.scala 11:37]
  wire [2:0] _T_1044 = _T_325 ? 3'h0 : _T_1043; // @[Lookup.scala 11:37]
  wire [2:0] _T_1045 = _T_321 ? 3'h0 : _T_1044; // @[Lookup.scala 11:37]
  wire [2:0] _T_1046 = _T_317 ? 3'h0 : _T_1045; // @[Lookup.scala 11:37]
  wire [2:0] _T_1047 = _T_313 ? 3'h0 : _T_1046; // @[Lookup.scala 11:37]
  wire [2:0] _T_1048 = _T_309 ? 3'h0 : _T_1047; // @[Lookup.scala 11:37]
  wire [2:0] _T_1049 = _T_305 ? 3'h0 : _T_1048; // @[Lookup.scala 11:37]
  wire [2:0] _T_1050 = _T_301 ? 3'h0 : _T_1049; // @[Lookup.scala 11:37]
  wire [2:0] _T_1051 = _T_297 ? 3'h0 : _T_1050; // @[Lookup.scala 11:37]
  wire [2:0] _T_1052 = _T_293 ? 3'h0 : _T_1051; // @[Lookup.scala 11:37]
  wire [2:0] _T_1053 = _T_289 ? 3'h0 : _T_1052; // @[Lookup.scala 11:37]
  wire [2:0] _T_1054 = _T_285 ? 3'h0 : _T_1053; // @[Lookup.scala 11:37]
  wire [2:0] _T_1055 = _T_281 ? 3'h0 : _T_1054; // @[Lookup.scala 11:37]
  wire [2:0] _T_1056 = _T_277 ? 3'h0 : _T_1055; // @[Lookup.scala 11:37]
  wire [2:0] _T_1057 = _T_273 ? 3'h0 : _T_1056; // @[Lookup.scala 11:37]
  wire [2:0] _T_1058 = _T_269 ? 3'h0 : _T_1057; // @[Lookup.scala 11:37]
  wire [2:0] _T_1059 = _T_265 ? 3'h0 : _T_1058; // @[Lookup.scala 11:37]
  wire [2:0] _T_1060 = _T_261 ? 3'h0 : _T_1059; // @[Lookup.scala 11:37]
  wire [2:0] _T_1061 = _T_257 ? 3'h0 : _T_1060; // @[Lookup.scala 11:37]
  wire [2:0] _T_1062 = _T_253 ? 3'h0 : _T_1061; // @[Lookup.scala 11:37]
  wire [2:0] _T_1063 = _T_249 ? 3'h0 : _T_1062; // @[Lookup.scala 11:37]
  wire [2:0] _T_1064 = _T_245 ? 3'h0 : _T_1063; // @[Lookup.scala 11:37]
  wire [2:0] _T_1065 = _T_241 ? 3'h0 : _T_1064; // @[Lookup.scala 11:37]
  wire [2:0] _T_1066 = _T_237 ? 3'h0 : _T_1065; // @[Lookup.scala 11:37]
  wire [2:0] cs0_6 = _T_233 ? 3'h0 : _T_1066; // @[Lookup.scala 11:37]
  wire  _T_1069 = _T_421 ? 1'h0 : _T_425; // @[Lookup.scala 11:37]
  wire  _T_1070 = _T_417 ? 1'h0 : _T_1069; // @[Lookup.scala 11:37]
  wire  _T_1071 = _T_413 ? 1'h0 : _T_1070; // @[Lookup.scala 11:37]
  wire  _T_1072 = _T_409 ? 1'h0 : _T_1071; // @[Lookup.scala 11:37]
  wire  _T_1073 = _T_405 ? 1'h0 : _T_1072; // @[Lookup.scala 11:37]
  wire  _T_1074 = _T_401 ? 1'h0 : _T_1073; // @[Lookup.scala 11:37]
  wire  _T_1075 = _T_397 ? 1'h0 : _T_1074; // @[Lookup.scala 11:37]
  wire  _T_1076 = _T_393 ? 1'h0 : _T_1075; // @[Lookup.scala 11:37]
  wire  _T_1077 = _T_389 ? 1'h0 : _T_1076; // @[Lookup.scala 11:37]
  wire  _T_1078 = _T_385 ? 1'h0 : _T_1077; // @[Lookup.scala 11:37]
  wire  _T_1079 = _T_381 ? 1'h0 : _T_1078; // @[Lookup.scala 11:37]
  wire  _T_1080 = _T_377 ? 1'h0 : _T_1079; // @[Lookup.scala 11:37]
  wire  _T_1081 = _T_373 ? 1'h0 : _T_1080; // @[Lookup.scala 11:37]
  wire  _T_1082 = _T_369 ? 1'h0 : _T_1081; // @[Lookup.scala 11:37]
  wire  _T_1083 = _T_365 ? 1'h0 : _T_1082; // @[Lookup.scala 11:37]
  wire  _T_1084 = _T_361 ? 1'h0 : _T_1083; // @[Lookup.scala 11:37]
  wire  _T_1085 = _T_357 ? 1'h0 : _T_1084; // @[Lookup.scala 11:37]
  wire  _T_1086 = _T_353 ? 1'h0 : _T_1085; // @[Lookup.scala 11:37]
  wire  _T_1087 = _T_349 ? 1'h0 : _T_1086; // @[Lookup.scala 11:37]
  wire  _T_1088 = _T_345 ? 1'h0 : _T_1087; // @[Lookup.scala 11:37]
  wire  _T_1089 = _T_341 ? 1'h0 : _T_1088; // @[Lookup.scala 11:37]
  wire  _T_1090 = _T_337 ? 1'h0 : _T_1089; // @[Lookup.scala 11:37]
  wire  _T_1091 = _T_333 ? 1'h0 : _T_1090; // @[Lookup.scala 11:37]
  wire  _T_1092 = _T_329 ? 1'h0 : _T_1091; // @[Lookup.scala 11:37]
  wire  _T_1093 = _T_325 ? 1'h0 : _T_1092; // @[Lookup.scala 11:37]
  wire  _T_1094 = _T_321 ? 1'h0 : _T_1093; // @[Lookup.scala 11:37]
  wire  _T_1095 = _T_317 ? 1'h0 : _T_1094; // @[Lookup.scala 11:37]
  wire  _T_1096 = _T_313 ? 1'h0 : _T_1095; // @[Lookup.scala 11:37]
  wire  _T_1097 = _T_309 ? 1'h0 : _T_1096; // @[Lookup.scala 11:37]
  wire  _T_1098 = _T_305 ? 1'h0 : _T_1097; // @[Lookup.scala 11:37]
  wire  _T_1099 = _T_301 ? 1'h0 : _T_1098; // @[Lookup.scala 11:37]
  wire  _T_1100 = _T_297 ? 1'h0 : _T_1099; // @[Lookup.scala 11:37]
  wire  _T_1101 = _T_293 ? 1'h0 : _T_1100; // @[Lookup.scala 11:37]
  wire  _T_1102 = _T_289 ? 1'h0 : _T_1101; // @[Lookup.scala 11:37]
  wire  _T_1103 = _T_285 ? 1'h0 : _T_1102; // @[Lookup.scala 11:37]
  wire  _T_1104 = _T_281 ? 1'h0 : _T_1103; // @[Lookup.scala 11:37]
  wire  _T_1105 = _T_277 ? 1'h0 : _T_1104; // @[Lookup.scala 11:37]
  wire  _T_1106 = _T_273 ? 1'h0 : _T_1105; // @[Lookup.scala 11:37]
  wire  _T_1107 = _T_269 ? 1'h0 : _T_1106; // @[Lookup.scala 11:37]
  wire  _T_1108 = _T_265 ? 1'h0 : _T_1107; // @[Lookup.scala 11:37]
  wire  _T_1109 = _T_261 ? 1'h0 : _T_1108; // @[Lookup.scala 11:37]
  wire  _T_1110 = _T_257 ? 1'h0 : _T_1109; // @[Lookup.scala 11:37]
  wire  _T_1111 = _T_253 ? 1'h0 : _T_1110; // @[Lookup.scala 11:37]
  wire  _T_1112 = _T_249 ? 1'h0 : _T_1111; // @[Lookup.scala 11:37]
  wire  _T_1113 = _T_245 ? 1'h0 : _T_1112; // @[Lookup.scala 11:37]
  wire  _T_1114 = _T_241 ? 1'h0 : _T_1113; // @[Lookup.scala 11:37]
  wire  _T_1115 = _T_237 ? 1'h0 : _T_1114; // @[Lookup.scala 11:37]
  wire  cs0_7 = _T_233 ? 1'h0 : _T_1115; // @[Lookup.scala 11:37]
  wire  _T_1116 = io_dat_exe_br_type == 4'h0; // @[cpath.scala 136:49]
  wire  _T_1117 = io_dat_exe_br_type == 4'h1; // @[cpath.scala 137:49]
  wire  _T_1119 = ~io_dat_exe_br_eq; // @[cpath.scala 137:65]
  wire [1:0] _T_1120 = _T_1119 ? 2'h1 : 2'h0; // @[cpath.scala 137:64]
  wire  _T_1121 = io_dat_exe_br_type == 4'h2; // @[cpath.scala 138:49]
  wire [1:0] _T_1122 = io_dat_exe_br_eq ? 2'h1 : 2'h0; // @[cpath.scala 138:64]
  wire  _T_1123 = io_dat_exe_br_type == 4'h3; // @[cpath.scala 139:49]
  wire  _T_1125 = ~io_dat_exe_br_lt; // @[cpath.scala 139:65]
  wire [1:0] _T_1126 = _T_1125 ? 2'h1 : 2'h0; // @[cpath.scala 139:64]
  wire  _T_1127 = io_dat_exe_br_type == 4'h4; // @[cpath.scala 140:49]
  wire  _T_1129 = ~io_dat_exe_br_ltu; // @[cpath.scala 140:65]
  wire [1:0] _T_1130 = _T_1129 ? 2'h1 : 2'h0; // @[cpath.scala 140:64]
  wire  _T_1131 = io_dat_exe_br_type == 4'h5; // @[cpath.scala 141:49]
  wire [1:0] _T_1132 = io_dat_exe_br_lt ? 2'h1 : 2'h0; // @[cpath.scala 141:64]
  wire  _T_1133 = io_dat_exe_br_type == 4'h6; // @[cpath.scala 142:49]
  wire [1:0] _T_1134 = io_dat_exe_br_ltu ? 2'h1 : 2'h0; // @[cpath.scala 142:64]
  wire  _T_1135 = io_dat_exe_br_type == 4'h7; // @[cpath.scala 143:49]
  wire  _T_1136 = io_dat_exe_br_type == 4'h8; // @[cpath.scala 144:49]
  wire [1:0] _T_1137 = _T_1136 ? 2'h2 : 2'h0; // @[cpath.scala 144:29]
  wire [1:0] _T_1138 = _T_1135 ? 2'h1 : _T_1137; // @[cpath.scala 143:29]
  wire [1:0] _T_1139 = _T_1133 ? _T_1134 : _T_1138; // @[cpath.scala 142:29]
  wire [1:0] _T_1140 = _T_1131 ? _T_1132 : _T_1139; // @[cpath.scala 141:29]
  wire [1:0] _T_1141 = _T_1127 ? _T_1130 : _T_1140; // @[cpath.scala 140:29]
  wire [1:0] _T_1142 = _T_1123 ? _T_1126 : _T_1141; // @[cpath.scala 139:29]
  wire [1:0] _T_1143 = _T_1121 ? _T_1122 : _T_1142; // @[cpath.scala 138:29]
  wire [1:0] _T_1144 = _T_1117 ? _T_1120 : _T_1143; // @[cpath.scala 137:29]
  wire [1:0] _T_1145 = _T_1116 ? 2'h0 : _T_1144; // @[cpath.scala 136:29]
  wire [1:0] ctrl_exe_pc_sel = io_ctl_pipeline_kill ? 2'h3 : _T_1145; // @[cpath.scala 135:29]
  wire  _T_1146 = ctrl_exe_pc_sel != 2'h0; // @[cpath.scala 148:35]
  wire  _T_1148 = ~io_imem_resp_valid; // @[cpath.scala 148:47]
  wire  _T_1149 = _T_1146 | _T_1148; // @[cpath.scala 148:44]
  wire  _T_1150 = _T_1149 | cs0_7; // @[cpath.scala 148:67]
  reg  _T_1152; // @[cpath.scala 148:86]
  wire  _T_1155 = ~cs_val_inst; // @[cpath.scala 155:25]
  wire  dec_exception = _T_1155 & io_imem_resp_valid; // @[cpath.scala 155:38]
  wire [4:0] dec_rs1_addr = io_dat_dec_inst[19:15]; // @[cpath.scala 160:38]
  wire [4:0] dec_rs2_addr = io_dat_dec_inst[24:20]; // @[cpath.scala 161:38]
  wire [4:0] dec_wbaddr = io_dat_dec_inst[11:7]; // @[cpath.scala 162:38]
  wire  dec_rs1_oen = _T_1146 ? 1'h0 : cs_rs1_oen; // @[cpath.scala 163:26]
  wire  dec_rs2_oen = _T_1146 ? 1'h0 : cs_rs2_oen; // @[cpath.scala 164:26]
  reg [4:0] exe_reg_wbaddr; // @[cpath.scala 166:33]
  reg  exe_reg_exception; // @[cpath.scala 172:33]
  reg  exe_reg_is_csr; // @[cpath.scala 174:28]
  reg  exe_inst_is_load; // @[cpath.scala 209:30]
  wire  _T_1198 = exe_reg_wbaddr == dec_rs1_addr; // @[cpath.scala 223:55]
  wire  _T_1199 = exe_inst_is_load & _T_1198; // @[cpath.scala 223:36]
  wire  _T_1201 = exe_reg_wbaddr != 5'h0; // @[cpath.scala 223:92]
  wire  _T_1202 = _T_1199 & _T_1201; // @[cpath.scala 223:73]
  wire  _T_1203 = _T_1202 & dec_rs1_oen; // @[cpath.scala 223:100]
  wire  _T_1204 = exe_reg_wbaddr == dec_rs2_addr; // @[cpath.scala 224:55]
  wire  _T_1205 = exe_inst_is_load & _T_1204; // @[cpath.scala 224:36]
  wire  _T_1208 = _T_1205 & _T_1201; // @[cpath.scala 224:73]
  wire  _T_1209 = _T_1208 & dec_rs2_oen; // @[cpath.scala 224:100]
  wire  _T_1210 = _T_1203 | _T_1209; // @[cpath.scala 223:116]
  wire  stall = _T_1210 | exe_reg_is_csr; // @[cpath.scala 224:116]
  wire  _T_1174 = ~stall; // @[cpath.scala 178:10]
  wire  _T_1214 = io_dat_mem_ctrl_dmem_val & io_dmem_resp_valid; // @[cpath.scala 244:53]
  wire  _T_1216 = ~io_dat_mem_ctrl_dmem_val; // @[cpath.scala 244:79]
  wire  _T_1217 = _T_1214 | _T_1216; // @[cpath.scala 244:76]
  wire  _T_1219 = ~_T_1217; // @[cpath.scala 244:41]
  wire  full_stall = _T_1148 | _T_1219; // @[cpath.scala 244:38]
  wire  _T_1176 = ~full_stall; // @[cpath.scala 178:20]
  wire  _T_1177 = _T_1174 & _T_1176; // @[cpath.scala 178:17]
  wire  _T_1182 = cs0_6 != 3'h0; // @[cpath.scala 191:44]
  wire  _T_1183 = cs0_6 != 3'h4; // @[cpath.scala 191:67]
  wire  _T_1184 = _T_1182 & _T_1183; // @[cpath.scala 191:53]
  wire  _T_1187 = stall & _T_1176; // @[cpath.scala 195:21]
  wire  _T_1196 = ~cs0_4; // @[cpath.scala 213:52]
  wire  _T_1197 = cs0_3 & _T_1196; // @[cpath.scala 213:37]
  reg  _T_1222; // @[cpath.scala 261:41]
  reg  _T_1225; // @[cpath.scala 263:31]
  wire  _T_1226 = cs0_6 == 3'h2; // @[cpath.scala 268:30]
  wire  _T_1227 = cs0_6 == 3'h3; // @[cpath.scala 268:54]
  wire  _T_1228 = _T_1226 | _T_1227; // @[cpath.scala 268:40]
  wire  _T_1230 = dec_rs1_addr == 5'h0; // @[cpath.scala 268:77]
  wire  csr_ren = _T_1228 & _T_1230; // @[cpath.scala 268:65]
  assign io_ctl_dec_stall = _T_1210 | exe_reg_is_csr; // @[cpath.scala 247:22]
  assign io_ctl_full_stall = _T_1148 | _T_1219; // @[cpath.scala 248:22]
  assign io_ctl_exe_pc_sel = io_ctl_pipeline_kill ? 2'h3 : _T_1145; // @[cpath.scala 249:22]
  assign io_ctl_br_type = _T_233 ? 4'h0 : _T_527; // @[cpath.scala 250:22]
  assign io_ctl_if_kill = _T_1150 | _T_1152; // @[cpath.scala 251:22]
  assign io_ctl_dec_kill = ctrl_exe_pc_sel != 2'h0; // @[cpath.scala 252:22]
  assign io_ctl_op1_sel = _T_233 ? 2'h0 : _T_576; // @[cpath.scala 253:22]
  assign io_ctl_op2_sel = _T_233 ? 3'h1 : _T_625; // @[cpath.scala 254:22]
  assign io_ctl_alu_fun = _T_233 ? 4'h0 : _T_772; // @[cpath.scala 255:22]
  assign io_ctl_wb_sel = _T_233 ? 2'h1 : _T_821; // @[cpath.scala 256:22]
  assign io_ctl_rf_wen = _T_233 | _T_870; // @[cpath.scala 257:22]
  assign io_ctl_mem_val = _T_233 | _T_919; // @[cpath.scala 274:22]
  assign io_ctl_mem_fcn = {{1'd0}, cs0_4}; // @[cpath.scala 275:22]
  assign io_ctl_mem_typ = _T_233 ? 3'h3 : _T_1017; // @[cpath.scala 276:21]
  assign io_ctl_csr_cmd = csr_ren ? 3'h5 : cs0_6; // @[cpath.scala 269:19]
  assign io_ctl_fencei = cs0_7 | _T_1222; // @[cpath.scala 261:22]
  assign io_ctl_pipeline_kill = io_dat_csr_eret | io_ctl_mem_exception; // @[cpath.scala 153:25]
  assign io_ctl_mem_exception = _T_1225; // @[cpath.scala 263:25]
  assign _GEN_111_0 = 32'h6013 == _T_232;
  assign _GEN_71_0 = 32'h1013 == _T_296;
  assign _GEN_324_0 = 32'h6013 == _T_232;
  assign _GEN_219_0 = 32'h37 == _T_264;
  assign _GEN_168_0 = 32'h5013 == _T_296;
  assign _GEN_1_0 = 32'h6063 == _T_232;
  assign _GEN_423_0 = reset;
  assign _GEN_44_0 = 32'h3 == _T_232;
  assign _GEN_267_0 = 32'h5013 == _T_296;
  assign _GEN_126_0 = 32'h67 == _T_232;
  assign _GEN_153_0 = 32'h5063 == _T_232;
  assign _GEN_225_0 = 32'h1003 == _T_232;
  assign _GEN_59_0 = 32'h5033 == _T_308;
  assign _GEN_252_0 = 32'h5063 == _T_232;
  assign _GEN_147_0 = 32'h1073 == _T_232;
  assign _GEN_351_0 = 32'h5063 == _T_232;
  assign _GEN_210_0 = 32'h5013 == _T_296;
  assign _GEN_246_0 = 32'h1073 == _T_232;
  assign _GEN_65_0 = 32'h2033 == _T_308;
  assign _GEN_132_0 = 32'h2013 == _T_232;
  assign _GEN_318_0 = 32'h5013 == _T_296;
  assign _GEN_92_0 = 32'h63 == _T_232;
  assign _GEN_345_0 = 32'h1073 == _T_232;
  assign _GEN_231_0 = 32'h5063 == _T_232;
  assign _GEN_417_0 = 32'h2003 == _T_232;
  assign _GEN_50_0 = 32'h5073 == _T_232;
  assign _GEN_330_0 = 32'h23 == _T_232;
  assign _GEN_86_0 = 32'h3 == _T_232;
  assign _GEN_339_0 = 32'h7b200073 == io_dat_dec_inst;
  assign _GEN_240_0 = 32'h7b200073 == io_dat_dec_inst;
  assign _GEN_234_0 = 32'h1023 == _T_232;
  assign _GEN_120_0 = 32'h1003 == _T_232;
  assign _GEN_129_0 = 32'h40005013 == _T_296;
  assign _GEN_333_0 = 32'h1003 == _T_232;
  assign _GEN_302_0 = 32'h7063 == _T_232;
  assign _GEN_228_0 = 32'h6063 == _T_232;
  assign _GEN_197_0 = 32'h63 == _T_232;
  assign _GEN_411_0 = ~full_stall;
  assign _GEN_401_0 = ctrl_exe_pc_sel != 2'h0;
  assign _GEN_47_0 = 32'h2073 == _T_232;
  assign _GEN_296_0 = 32'h2073 == _T_232;
  assign _GEN_74_0 = 32'h4013 == _T_232;
  assign _GEN_213_0 = 32'h3013 == _T_232;
  assign _GEN_32_0 = 32'h4013 == _T_232;
  assign _GEN_68_0 = 32'h1033 == _T_308;
  assign _GEN_135_0 = 32'h7013 == _T_232;
  assign _GEN_26_0 = 32'h1033 == _T_308;
  assign _GEN_53_0 = 32'h7063 == _T_232;
  assign _GEN_141_0 = 32'h4003 == _T_232;
  assign _GEN_327_0 = 32'h37 == _T_264;
  assign _GEN_395_0 = io_dat_exe_br_type == 4'h4;
  assign _GEN_249_0 = 32'h6063 == _T_232;
  assign _GEN_114_0 = 32'h37 == _T_264;
  assign _GEN_312_0 = 32'h7033 == _T_308;
  assign _GEN_203_0 = 32'h6033 == _T_308;
  assign _GEN_20_0 = 32'h6033 == _T_308;
  assign _GEN_15_0 = 32'h67 == _T_232;
  assign _GEN_216_0 = 32'h6013 == _T_232;
  assign _GEN_206_0 = 32'h2033 == _T_308;
  assign _GEN_420_0 = 32'h2003 == _T_232;
  assign _GEN_123_0 = 32'h6f == _T_264;
  assign _GEN_315_0 = 32'h40000033 == _T_308;
  assign _GEN_284_0 = 32'h23 == _T_232;
  assign _GEN_179_0 = 32'h1023 == _T_232;
  assign _GEN_222_0 = 32'h23 == _T_232;
  assign _GEN_377_0 = 32'h1023 == _T_232;
  assign _GEN_191_0 = 32'h5073 == _T_232;
  assign _GEN_290_0 = 32'h100073 == io_dat_dec_inst;
  assign _GEN_404_0 = ctrl_exe_pc_sel != 2'h0;
  assign _GEN_56_1 = 32'h63 == _T_232;
  assign _GEN_305_0 = 32'h63 == _T_232;
  assign _GEN_299_0 = 32'h5073 == _T_232;
  assign _GEN_185_0 = 32'h3 == _T_232;
  assign _GEN_398_0 = io_dat_exe_br_type == 4'h1;
  assign _GEN_41_0 = 32'h5003 == _T_232;
  assign _GEN_321_0 = 32'h3013 == _T_232;
  assign _GEN_414_0 = 32'h2003 == _T_232;
  assign _GEN_383_0 = 32'h3 == _T_232;
  assign _GEN_35_0 = 32'h13 == _T_232;
  assign _GEN_29_0 = 32'h1013 == _T_296;
  assign _GEN_278_0 = 32'h5003 == _T_232;
  assign _GEN_117_0 = 32'h23 == _T_232;
  assign _GEN_365_0 = 32'h1033 == _T_308;
  assign _GEN_359_0 = 32'h6033 == _T_308;
  assign _GEN_38_0 = 32'h1023 == _T_232;
  assign _GEN_167_0 = 32'h1033 == _T_308;
  assign _GEN_350_0 = 32'h7063 == _T_232;
  assign _GEN_106_0 = 32'h40005013 == _T_296;
  assign _GEN_18_0 = 32'h40005033 == _T_308;
  assign _GEN_293_0 = 32'h73 == io_dat_dec_inst;
  assign _GEN_371_0 = 32'h4013 == _T_232;
  assign _GEN_251_0 = 32'h7063 == _T_232;
  assign _GEN_209_0 = 32'h1033 == _T_308;
  assign _GEN_308_0 = 32'h5033 == _T_308;
  assign _GEN_173_0 = 32'h4013 == _T_232;
  assign _GEN_200_0 = 32'h5033 == _T_308;
  assign _GEN_386_0 = io_dat_exe_br_eq;
  assign _GEN_272_0 = 32'h4013 == _T_232;
  assign _GEN_91_1 = 32'h1063 == _T_232;
  assign _GEN_194_0 = 32'h7063 == _T_232;
  assign _GEN_188_0 = 32'h2073 == _T_232;
  assign _GEN_392_0 = io_dat_exe_br_type == 4'h7;
  assign _GEN_23_0 = 32'h2033 == _T_308;
  assign _GEN_407_0 = stall & _T_1176;
  assign _GEN_287_0 = 32'h1003 == _T_232;
  assign _GEN_266_0 = 32'h1033 == _T_308;
  assign _GEN_374_0 = 32'h13 == _T_232;
  assign _GEN_233_0 = 32'h63 == _T_232;
  assign _GEN_269_0 = 32'h1013 == _T_296;
  assign _GEN_260_0 = 32'h6033 == _T_308;
  assign _GEN_161_0 = 32'h6033 == _T_308;
  assign _GEN_155_0 = 32'h63 == _T_232;
  assign _GEN_368_0 = 32'h1013 == _T_296;
  assign _GEN_254_0 = 32'h63 == _T_232;
  assign _GEN_281_0 = 32'h3 == _T_232;
  assign _GEN_73_0 = 32'h2013 == _T_232;
  assign _GEN_353_0 = 32'h63 == _T_232;
  assign _GEN_332_0 = 32'h5003 == _T_232;
  assign _GEN_88_1 = 32'h4063 == _T_232;
  assign _GEN_176_0 = 32'h13 == _T_232;
  assign _GEN_380_0 = 32'h5003 == _T_232;
  assign _GEN_389_0 = io_dat_exe_br_lt;
  assign _GEN_94_0 = 32'h6f == _T_264;
  assign _GEN_347_0 = 32'h5073 == _T_232;
  assign _GEN_109_0 = 32'h2013 == _T_232;
  assign _GEN_182_0 = 32'h5003 == _T_232;
  assign _GEN_9_0 = 32'h5063 == _T_232;
  assign _GEN_149_0 = 32'h5073 == _T_232;
  assign _GEN_248_0 = 32'h5073 == _T_232;
  assign _GEN_275_0 = 32'h13 == _T_232;
  assign _GEN_140_1 = 32'h1003 == _T_232;
  assign _GEN_100_0 = 32'h3033 == _T_308;
  assign _GEN_362_0 = 32'h2033 == _T_308;
  assign _GEN_413_0 = 32'h2003 == _T_232;
  assign _GEN_76_0 = 32'h7013 == _T_232;
  assign _GEN_164_0 = 32'h2033 == _T_308;
  assign _GEN_242_0 = 32'h73 == io_dat_dec_inst;
  assign _GEN_137_0 = 32'h37 == _T_264;
  assign _GEN_341_0 = 32'h73 == io_dat_dec_inst;
  assign _GEN_263_0 = 32'h2033 == _T_308;
  assign _GEN_257_0 = 32'h5033 == _T_308;
  assign _GEN_122_1 = 32'h3 == _T_232;
  assign _GEN_143_0 = 32'h2003 == _T_232;
  assign _GEN_82_0 = 32'h2023 == _T_232;
  assign _GEN_170_0 = 32'h1013 == _T_296;
  assign _GEN_356_0 = 32'h5033 == _T_308;
  assign _GEN_221_0 = 32'h1023 == _T_232;
  assign _GEN_215_0 = 32'h4013 == _T_232;
  assign _GEN_320_0 = 32'h1013 == _T_296;
  assign _GEN_314_0 = 32'h2033 == _T_308;
  assign _GEN_329_0 = 32'h1023 == _T_232;
  assign _GEN_103_1 = 32'h33 == _T_308;
  assign _GEN_97_0 = 32'h4033 == _T_308;
  assign _GEN_236_0 = 32'h2023 == _T_232;
  assign _GEN_61_0 = 32'h4033 == _T_308;
  assign _GEN_55_0 = 32'h1063 == _T_232;
  assign _GEN_335_0 = 32'h3 == _T_232;
  assign _GEN_158_0 = 32'h5033 == _T_308;
  assign _GEN_422_0 = reset;
  assign _GEN_245_0 = 32'h2073 == _T_232;
  assign _GEN_37_0 = 32'h17 == _T_264;
  assign _GEN_125_1 = 32'h17 == _T_264;
  assign _GEN_70_0 = 32'h40005013 == _T_296;
  assign _GEN_64_0 = 32'h3033 == _T_308;
  assign _GEN_344_0 = 32'h2073 == _T_232;
  assign _GEN_338_0 = 32'h100073 == io_dat_dec_inst;
  assign _GEN_416_0 = 32'h2003 == _T_232;
  assign _GEN_406_1 = stall & _T_1176;
  assign _GEN_58_0 = 32'h6f == _T_264;
  assign _GEN_85_1 = 32'h4003 == _T_232;
  assign _GEN_43_0 = 32'h4003 == _T_232;
  assign _GEN_131_0 = 32'h3013 == _T_232;
  assign _GEN_230_0 = 32'h7063 == _T_232;
  assign _GEN_239_0 = 32'h100073 == io_dat_dec_inst;
  assign _GEN_152_0 = 32'h7063 == _T_232;
  assign _GEN_307_1 = 32'h6f == _T_264;
  assign _GEN_146_1 = 32'h2073 == _T_232;
  assign _GEN_224_0 = 32'h5003 == _T_232;
  assign _GEN_110_0 = 32'h4013 == _T_232;
  assign _GEN_119_1 = 32'h5003 == _T_232;
  assign _GEN_323_0 = 32'h4013 == _T_232;
  assign _GEN_317_0 = 32'h1033 == _T_308;
  assign _GEN_79_1 = 32'h17 == _T_264;
  assign _GEN_218_0 = 32'h13 == _T_232;
  assign _GEN_208_0 = 32'h33 == _T_308;
  assign _GEN_196_0 = 32'h1063 == _T_232;
  assign _GEN_31_0 = 32'h2013 == _T_232;
  assign _GEN_400_0 = io_ctl_pipeline_kill;
  assign _GEN_113_1 = 32'h13 == _T_232;
  assign _GEN_212_0 = 32'h1013 == _T_296;
  assign _GEN_181_0 = 32'h2023 == _T_232;
  assign _GEN_227_0 = 32'h3 == _T_232;
  assign _GEN_425_0 = 32'h2003 == _T_232;
  assign _GEN_280_0 = 32'h4003 == _T_232;
  assign _GEN_46_0 = 32'h3073 == _T_232;
  assign _GEN_134_0 = 32'h6013 == _T_232;
  assign _GEN_289_0 = 32'h3 == _T_232;
  assign _GEN_202_0 = 32'h4033 == _T_308;
  assign _GEN_419_0 = _T_1228 & _T_1230;
  assign _GEN_388_0 = ~io_dat_exe_br_ltu;
  assign _GEN_410_0 = _T_1174 & _T_1176;
  assign _GEN_52_0 = 32'h4063 == _T_232;
  assign _GEN_311_0 = 32'h6033 == _T_308;
  assign _GEN_301_0 = 32'h4063 == _T_232;
  assign _GEN_295_0 = 32'h3073 == _T_232;
  assign _GEN_67_0 = 32'h33 == _T_308;
  assign _GEN_25_0 = 32'h33 == _T_308;
  assign _GEN_409_1 = _T_1174 & _T_1176;
  assign _GEN_326_0 = 32'h13 == _T_232;
  assign _GEN_394_0 = io_dat_exe_br_type == 4'h5;
  assign _GEN_128_0 = 32'h5013 == _T_296;
  assign _GEN_376_0 = 32'h17 == _T_264;
  assign _GEN_40_0 = 32'h2023 == _T_232;
  assign _GEN_34_0 = 32'h7013 == _T_232;
  assign _GEN_49_0 = 32'h6073 == _T_232;
  assign _GEN_102_0 = 32'h40000033 == _T_308;
  assign _GEN_190_0 = 32'h6073 == _T_232;
  assign _GEN_205_0 = 32'h3033 == _T_308;
  assign _GEN_298_0 = 32'h6073 == _T_232;
  assign _GEN_163_1 = 32'h3033 == _T_308;
  assign _GEN_14_0 = 32'h63 == _T_232;
  assign _GEN_116_0 = 32'h1023 == _T_232;
  assign _GEN_283_0 = 32'h1023 == _T_232;
  assign _GEN_184_0 = 32'h4003 == _T_232;
  assign _GEN_178_1 = 32'h17 == _T_264;
  assign _GEN_382_0 = 32'h4003 == _T_232;
  assign _GEN_397_0 = io_dat_exe_br_type == 4'h2;
  assign _GEN_277_0 = 32'h17 == _T_264;
  assign _GEN_304_1 = 32'h1063 == _T_232;
  assign _GEN_199_0 = 32'h6f == _T_264;
  assign _GEN_403_0 = ctrl_exe_pc_sel != 2'h0;
  assign _GEN_262_0 = 32'h3033 == _T_308;
  assign _GEN_28_0 = 32'h40005013 == _T_296;
  assign _GEN_361_0 = 32'h3033 == _T_308;
  assign _GEN_96_0 = 32'h40005033 == _T_308;
  assign _GEN_193_0 = 32'h4063 == _T_232;
  assign _GEN_379_0 = 32'h2023 == _T_232;
  assign _GEN_244_1 = 32'h3073 == _T_232;
  assign _GEN_271_0 = 32'h2013 == _T_232;
  assign _GEN_151_2 = 32'h4063 == _T_232;
  assign _GEN_166_1 = 32'h33 == _T_308;
  assign _GEN_370_0 = 32'h2013 == _T_232;
  assign _GEN_364_0 = 32'h33 == _T_308;
  assign _GEN_259_0 = 32'h4033 == _T_308;
  assign _GEN_292_0 = 32'h30200073 == io_dat_dec_inst;
  assign _GEN_84_0 = 32'h1003 == _T_232;
  assign _GEN_78_0 = 32'h37 == _T_264;
  assign _GEN_385_0 = ~io_dat_exe_br_eq;
  assign _GEN_250_0 = 32'h4063 == _T_232;
  assign _GEN_343_0 = 32'h3073 == _T_232;
  assign _GEN_105_0 = 32'h5013 == _T_296;
  assign _GEN_99_0 = 32'h7033 == _T_308;
  assign _GEN_358_0 = 32'h4033 == _T_308;
  assign _GEN_22_0 = 32'h3033 == _T_308;
  assign _GEN_265_0 = 32'h33 == _T_308;
  assign _GEN_17_0 = 32'h5033 == _T_308;
  assign _GEN_90_1 = 32'h5063 == _T_232;
  assign _GEN_172_1 = 32'h2013 == _T_232;
  assign _GEN_187_0 = 32'h3073 == _T_232;
  assign _GEN_391_0 = io_dat_exe_br_type == 4'h8;
  assign _GEN_286_0 = 32'h5003 == _T_232;
  assign _GEN_145_1 = 32'h3073 == _T_232;
  assign _GEN_232_0 = 32'h1063 == _T_232;
  assign _GEN_274_0 = 32'h7013 == _T_232;
  assign _GEN_175_1 = 32'h7013 == _T_232;
  assign _GEN_169_1 = 32'h40005013 == _T_296;
  assign _GEN_247_0 = 32'h6073 == _T_232;
  assign _GEN_133_1 = 32'h4013 == _T_232;
  assign _GEN_160_1 = 32'h4033 == _T_308;
  assign _GEN_346_0 = 32'h6073 == _T_232;
  assign _GEN_373_0 = 32'h7013 == _T_232;
  assign _GEN_424_1 = reset;
  assign _GEN_268_0 = 32'h40005013 == _T_296;
  assign _GEN_127_1 = 32'h6f == _T_264;
  assign _GEN_8_0 = 32'h7063 == _T_232;
  assign _GEN_331_1 = 32'h2023 == _T_232;
  assign _GEN_93_1 = 32'h67 == _T_232;
  assign _GEN_87_1 = 32'h6063 == _T_232;
  assign _GEN_367_0 = 32'h40005013 == _T_296;
  assign _GEN_226_0 = 32'h4003 == _T_232;
  assign _GEN_253_1 = 32'h1063 == _T_232;
  assign _GEN_325_1 = 32'h7013 == _T_232;
  assign _GEN_148_1 = 32'h6073 == _T_232;
  assign _GEN_352_1 = 32'h1063 == _T_232;
  assign _GEN_108_0 = 32'h3013 == _T_232;
  assign _GEN_72_1 = 32'h3013 == _T_232;
  assign _GEN_66_0 = 32'h40000033 == _T_308;
  assign _GEN_154_1 = 32'h1063 == _T_232;
  assign _GEN_241_0 = 32'h30200073 == io_dat_dec_inst;
  assign _GEN_402_1 = ctrl_exe_pc_sel != 2'h0;
  assign _GEN_48_0 = 32'h1073 == _T_232;
  assign _GEN_60_0 = 32'h40005033 == _T_308;
  assign _GEN_75_1 = 32'h6013 == _T_232;
  assign _GEN_349_0 = 32'h4063 == _T_232;
  assign _GEN_214_0 = 32'h2013 == _T_232;
  assign _GEN_412_1 = io_ctl_pipeline_kill;
  assign _GEN_256_0 = 32'h6f == _T_264;
  assign _GEN_121_1 = 32'h4003 == _T_232;
  assign _GEN_81_0 = 32'h23 == _T_232;
  assign _GEN_54_0 = 32'h5063 == _T_232;
  assign _GEN_136_1 = 32'h13 == _T_232;
  assign _GEN_142_1 = 32'h3 == _T_232;
  assign _GEN_340_0 = 32'h30200073 == io_dat_dec_inst;
  assign _GEN_355_0 = 32'h6f == _T_264;
  assign _GEN_235_0 = 32'h23 == _T_232;
  assign _GEN_313_1 = 32'h3033 == _T_308;
  assign _GEN_69_1 = 32'h5013 == _T_296;
  assign _GEN_157_1 = 32'h6f == _T_264;
  assign _GEN_220_0 = 32'h17 == _T_264;
  assign _GEN_229_0 = 32'h4063 == _T_232;
  assign _GEN_115_1 = 32'h17 == _T_264;
  assign _GEN_334_0 = 32'h4003 == _T_232;
  assign _GEN_328_0 = 32'h17 == _T_264;
  assign _GEN_36_0 = 32'h37 == _T_264;
  assign _GEN_405_1 = ctrl_exe_pc_sel != 2'h0;
  assign _GEN_415_1 = 32'h2003 == _T_232;
  assign _GEN_124_1 = 32'h37 == _T_264;
  assign _GEN_322_0 = 32'h2013 == _T_232;
  assign _GEN_337_1 = 32'h10500073 == io_dat_dec_inst;
  assign _GEN_223_0 = 32'h2023 == _T_232;
  assign _GEN_217_0 = 32'h7013 == _T_232;
  assign _GEN_192_0 = 32'h6063 == _T_232;
  assign _GEN_390_1 = io_dat_exe_br_ltu;
  assign _GEN_42_1 = 32'h1003 == _T_232;
  assign _GEN_291_1 = 32'h7b200073 == io_dat_dec_inst;
  assign _GEN_139_1 = 32'h5003 == _T_232;
  assign _GEN_207_0 = 32'h40000033 == _T_308;
  assign _GEN_399_1 = io_dat_exe_br_type == 4'h0;
  assign _GEN_421_0 = _T_1174 & _T_1176;
  assign _GEN_63_0 = 32'h7033 == _T_308;
  assign _GEN_316_1 = 32'h33 == _T_308;
  assign _GEN_306_1 = 32'h67 == _T_232;
  assign _GEN_21_1 = 32'h7033 == _T_308;
  assign _GEN_384_1 = 32'h2003 == _T_232;
  assign _GEN_118_1 = 32'h2023 == _T_232;
  assign _GEN_57_0 = 32'h67 == _T_232;
  assign _GEN_130_1 = 32'h1013 == _T_296;
  assign _GEN_238_1 = 32'h10500073 == io_dat_dec_inst;
  assign _GEN_45_1 = 32'h7073 == _T_232;
  assign _GEN_201_0 = 32'h40005033 == _T_308;
  assign _GEN_195_0 = 32'h5063 == _T_232;
  assign _GEN_309_1 = 32'h40005033 == _T_308;
  assign _GEN_372_1 = 32'h6013 == _T_232;
  assign _GEN_19_0 = 32'h4033 == _T_308;
  assign _GEN_51_0 = 32'h6063 == _T_232;
  assign _GEN_294_1 = 32'h7073 == _T_232;
  assign _GEN_180_0 = 32'h23 == _T_232;
  assign _GEN_189_0 = 32'h1073 == _T_232;
  assign _GEN_211_0 = 32'h40005013 == _T_296;
  assign _GEN_393_1 = io_dat_exe_br_type == 4'h6;
  assign _GEN_387_1 = ~io_dat_exe_br_lt;
  assign _GEN_39_0 = 32'h23 == _T_232;
  assign _GEN_288_1 = 32'h4003 == _T_232;
  assign _GEN_310_1 = 32'h4033 == _T_308;
  assign _GEN_300_1 = 32'h6063 == _T_232;
  assign _GEN_319_1 = 32'h40005013 == _T_296;
  assign _GEN_107_1 = 32'h1013 == _T_296;
  assign _GEN_174_1 = 32'h6013 == _T_232;
  assign _GEN_30_0 = 32'h3013 == _T_232;
  assign _GEN_24_0 = 32'h40000033 == _T_308;
  assign _GEN_408_1 = stall & _T_1176;
  assign _GEN_418_1 = 32'h2003 == _T_232;
  assign _GEN_273_1 = 32'h6013 == _T_232;
  assign _GEN_5_1 = 32'h4063 == _T_232;
  assign _GEN_112_1 = 32'h7013 == _T_232;
  assign _GEN_366_1 = 32'h5013 == _T_296;
  assign _GEN_360_1 = 32'h7033 == _T_308;
  assign _GEN_354_1 = 32'h67 == _T_232;
  assign _GEN_33_1 = 32'h6013 == _T_232;
  assign _GEN_276_1 = 32'h37 == _T_264;
  assign _GEN_348_1 = 32'h6063 == _T_232;
  assign _GEN_101_1 = 32'h2033 == _T_308;
  assign _GEN_375_1 = 32'h37 == _T_264;
  assign _GEN_27_0 = 32'h5013 == _T_296;
  assign _GEN_13_0 = 32'h1063 == _T_232;
  assign _GEN_297_1 = 32'h1073 == _T_232;
  assign _GEN_89_1 = 32'h7063 == _T_232;
  assign _GEN_177_1 = 32'h37 == _T_264;
  assign _GEN_255_1 = 32'h67 == _T_232;
  assign _GEN_204_0 = 32'h7033 == _T_308;
  assign _GEN_80_1 = 32'h1023 == _T_232;
  assign _GEN_303_1 = 32'h5063 == _T_232;
  assign _GEN_162_1 = 32'h7033 == _T_308;
  assign _GEN_198_0 = 32'h67 == _T_232;
  assign _GEN_381_1 = 32'h1003 == _T_232;
  assign _GEN_261_1 = 32'h7033 == _T_308;
  assign _GEN_156_1 = 32'h67 == _T_232;
  assign _GEN_95_1 = 32'h5033 == _T_308;
  assign _GEN_183_0 = 32'h1003 == _T_232;
  assign _GEN_369_1 = 32'h3013 == _T_232;
  assign _GEN_282_1 = 32'h2003 == _T_232;
  assign _GEN_396_1 = io_dat_exe_br_type == 4'h3;
  assign _GEN_378_1 = 32'h23 == _T_232;
  assign _GEN_186_0 = 32'h7073 == _T_232;
  assign _GEN_62_0 = 32'h6033 == _T_308;
  assign _GEN_285_1 = 32'h2023 == _T_232;
  assign _GEN_336_1 = 32'h2003 == _T_232;
  assign _GEN_144_1 = 32'h7073 == _T_232;
  assign _GEN_150_2 = 32'h6063 == _T_232;
  assign _GEN_363_1 = 32'h40000033 == _T_308;
  assign _GEN_243_1 = 32'h7073 == _T_232;
  assign _GEN_258_1 = 32'h40005033 == _T_308;
  assign _GEN_138_1 = 32'h17 == _T_264;
  assign _GEN_171_1 = 32'h3013 == _T_232;
  assign _GEN_357_1 = 32'h40005033 == _T_308;
  assign _GEN_165_1 = 32'h40000033 == _T_308;
  assign _GEN_264_1 = 32'h40000033 == _T_308;
  assign _GEN_16_1 = 32'h6f == _T_264;
  assign _GEN_342_1 = 32'h7073 == _T_232;
  assign _GEN_98_1 = 32'h6033 == _T_308;
  assign _GEN_237_1 = 32'h100f == _T_232;
  assign _GEN_83_1 = 32'h5003 == _T_232;
  assign _GEN_77_0 = 32'h13 == _T_232;
  assign _GEN_270_1 = 32'h3013 == _T_232;
  assign _GEN_279_1 = 32'h1003 == _T_232;
  assign _GEN_159_1 = 32'h40005033 == _T_308;
  assign _GEN_104_1 = 32'h1033 == _T_308;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1152 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  exe_reg_wbaddr = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  exe_reg_exception = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  exe_reg_is_csr = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  exe_inst_is_load = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_1222 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_1225 = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_1152 <= 1'h0;
    end else if (_T_233) begin
      _T_1152 <= 1'h0;
    end else if (_T_237) begin
      _T_1152 <= 1'h0;
    end else if (_T_241) begin
      _T_1152 <= 1'h0;
    end else if (_T_245) begin
      _T_1152 <= 1'h0;
    end else if (_T_249) begin
      _T_1152 <= 1'h0;
    end else if (_T_253) begin
      _T_1152 <= 1'h0;
    end else if (_T_257) begin
      _T_1152 <= 1'h0;
    end else if (_T_261) begin
      _T_1152 <= 1'h0;
    end else if (_T_265) begin
      _T_1152 <= 1'h0;
    end else if (_T_269) begin
      _T_1152 <= 1'h0;
    end else if (_T_273) begin
      _T_1152 <= 1'h0;
    end else if (_T_277) begin
      _T_1152 <= 1'h0;
    end else if (_T_281) begin
      _T_1152 <= 1'h0;
    end else if (_T_285) begin
      _T_1152 <= 1'h0;
    end else if (_T_289) begin
      _T_1152 <= 1'h0;
    end else if (_T_293) begin
      _T_1152 <= 1'h0;
    end else if (_T_297) begin
      _T_1152 <= 1'h0;
    end else if (_T_301) begin
      _T_1152 <= 1'h0;
    end else if (_T_305) begin
      _T_1152 <= 1'h0;
    end else if (_T_309) begin
      _T_1152 <= 1'h0;
    end else if (_T_313) begin
      _T_1152 <= 1'h0;
    end else if (_T_317) begin
      _T_1152 <= 1'h0;
    end else if (_T_321) begin
      _T_1152 <= 1'h0;
    end else if (_T_325) begin
      _T_1152 <= 1'h0;
    end else if (_T_329) begin
      _T_1152 <= 1'h0;
    end else if (_T_333) begin
      _T_1152 <= 1'h0;
    end else if (_T_337) begin
      _T_1152 <= 1'h0;
    end else if (_T_341) begin
      _T_1152 <= 1'h0;
    end else if (_T_345) begin
      _T_1152 <= 1'h0;
    end else if (_T_349) begin
      _T_1152 <= 1'h0;
    end else if (_T_353) begin
      _T_1152 <= 1'h0;
    end else if (_T_357) begin
      _T_1152 <= 1'h0;
    end else if (_T_361) begin
      _T_1152 <= 1'h0;
    end else if (_T_365) begin
      _T_1152 <= 1'h0;
    end else if (_T_369) begin
      _T_1152 <= 1'h0;
    end else if (_T_373) begin
      _T_1152 <= 1'h0;
    end else if (_T_377) begin
      _T_1152 <= 1'h0;
    end else if (_T_381) begin
      _T_1152 <= 1'h0;
    end else if (_T_385) begin
      _T_1152 <= 1'h0;
    end else if (_T_389) begin
      _T_1152 <= 1'h0;
    end else if (_T_393) begin
      _T_1152 <= 1'h0;
    end else if (_T_397) begin
      _T_1152 <= 1'h0;
    end else if (_T_401) begin
      _T_1152 <= 1'h0;
    end else if (_T_405) begin
      _T_1152 <= 1'h0;
    end else if (_T_409) begin
      _T_1152 <= 1'h0;
    end else if (_T_413) begin
      _T_1152 <= 1'h0;
    end else if (_T_417) begin
      _T_1152 <= 1'h0;
    end else if (_T_421) begin
      _T_1152 <= 1'h0;
    end else begin
      _T_1152 <= _T_425;
    end
    if (metaReset) begin
      exe_reg_wbaddr <= 5'h0;
    end else if (_T_1177) begin
      if (_T_1146) begin
        exe_reg_wbaddr <= 5'h0;
      end else begin
        exe_reg_wbaddr <= dec_wbaddr;
      end
    end else if (_T_1187) begin
      exe_reg_wbaddr <= 5'h0;
    end
    if (metaReset) begin
      exe_reg_exception <= 1'h0;
    end else if (reset) begin
      exe_reg_exception <= 1'h0;
    end else if (_T_1177) begin
      if (_T_1146) begin
        exe_reg_exception <= 1'h0;
      end else begin
        exe_reg_exception <= dec_exception;
      end
    end else if (_T_1187) begin
      exe_reg_exception <= 1'h0;
    end
    if (metaReset) begin
      exe_reg_is_csr <= 1'h0;
    end else if (reset) begin
      exe_reg_is_csr <= 1'h0;
    end else if (_T_1177) begin
      if (_T_1146) begin
        exe_reg_is_csr <= 1'h0;
      end else begin
        exe_reg_is_csr <= _T_1184;
      end
    end else if (_T_1187) begin
      exe_reg_is_csr <= 1'h0;
    end
    if (metaReset) begin
      exe_inst_is_load <= 1'h0;
    end else if (reset) begin
      exe_inst_is_load <= 1'h0;
    end else if (_T_1176) begin
      exe_inst_is_load <= _T_1197;
    end
    if (metaReset) begin
      _T_1222 <= 1'h0;
    end else if (_T_233) begin
      _T_1222 <= 1'h0;
    end else if (_T_237) begin
      _T_1222 <= 1'h0;
    end else if (_T_241) begin
      _T_1222 <= 1'h0;
    end else if (_T_245) begin
      _T_1222 <= 1'h0;
    end else if (_T_249) begin
      _T_1222 <= 1'h0;
    end else if (_T_253) begin
      _T_1222 <= 1'h0;
    end else if (_T_257) begin
      _T_1222 <= 1'h0;
    end else if (_T_261) begin
      _T_1222 <= 1'h0;
    end else if (_T_265) begin
      _T_1222 <= 1'h0;
    end else if (_T_269) begin
      _T_1222 <= 1'h0;
    end else if (_T_273) begin
      _T_1222 <= 1'h0;
    end else if (_T_277) begin
      _T_1222 <= 1'h0;
    end else if (_T_281) begin
      _T_1222 <= 1'h0;
    end else if (_T_285) begin
      _T_1222 <= 1'h0;
    end else if (_T_289) begin
      _T_1222 <= 1'h0;
    end else if (_T_293) begin
      _T_1222 <= 1'h0;
    end else if (_T_297) begin
      _T_1222 <= 1'h0;
    end else if (_T_301) begin
      _T_1222 <= 1'h0;
    end else if (_T_305) begin
      _T_1222 <= 1'h0;
    end else if (_T_309) begin
      _T_1222 <= 1'h0;
    end else if (_T_313) begin
      _T_1222 <= 1'h0;
    end else if (_T_317) begin
      _T_1222 <= 1'h0;
    end else if (_T_321) begin
      _T_1222 <= 1'h0;
    end else if (_T_325) begin
      _T_1222 <= 1'h0;
    end else if (_T_329) begin
      _T_1222 <= 1'h0;
    end else if (_T_333) begin
      _T_1222 <= 1'h0;
    end else if (_T_337) begin
      _T_1222 <= 1'h0;
    end else if (_T_341) begin
      _T_1222 <= 1'h0;
    end else if (_T_345) begin
      _T_1222 <= 1'h0;
    end else if (_T_349) begin
      _T_1222 <= 1'h0;
    end else if (_T_353) begin
      _T_1222 <= 1'h0;
    end else if (_T_357) begin
      _T_1222 <= 1'h0;
    end else if (_T_361) begin
      _T_1222 <= 1'h0;
    end else if (_T_365) begin
      _T_1222 <= 1'h0;
    end else if (_T_369) begin
      _T_1222 <= 1'h0;
    end else if (_T_373) begin
      _T_1222 <= 1'h0;
    end else if (_T_377) begin
      _T_1222 <= 1'h0;
    end else if (_T_381) begin
      _T_1222 <= 1'h0;
    end else if (_T_385) begin
      _T_1222 <= 1'h0;
    end else if (_T_389) begin
      _T_1222 <= 1'h0;
    end else if (_T_393) begin
      _T_1222 <= 1'h0;
    end else if (_T_397) begin
      _T_1222 <= 1'h0;
    end else if (_T_401) begin
      _T_1222 <= 1'h0;
    end else if (_T_405) begin
      _T_1222 <= 1'h0;
    end else if (_T_409) begin
      _T_1222 <= 1'h0;
    end else if (_T_413) begin
      _T_1222 <= 1'h0;
    end else if (_T_417) begin
      _T_1222 <= 1'h0;
    end else if (_T_421) begin
      _T_1222 <= 1'h0;
    end else begin
      _T_1222 <= _T_425;
    end
    if (metaReset) begin
      _T_1225 <= 1'h0;
    end else begin
      _T_1225 <= exe_reg_exception;
    end
  end
endmodule
module RegisterFile(
  input         metaReset,
  input         clock,
  input  [4:0]  io_rs1_addr,
  output [31:0] io_rs1_data,
  input  [4:0]  io_rs2_addr,
  output [31:0] io_rs2_data,
  input  [4:0]  io_waddr,
  input  [31:0] io_wdata,
  input         io_wen,
  output        _GEN_0_0,
  output        _GEN_1_3
);
  wire  mem_sparse_metaReset;
  wire  mem_sparse_clock;
  wire [4:0] mem_sparse_io_w_0_addr;
  wire  mem_sparse_io_w_0_en;
  wire [31:0] mem_sparse_io_w_0_data;
  wire [4:0] mem_sparse_io_r_0_addr;
  wire [31:0] mem_sparse_io_r_0_data;
  wire [4:0] mem_sparse_io_r_1_addr;
  wire [31:0] mem_sparse_io_r_1_data;
  wire  _T_18 = io_waddr != 5'h0; // @[regfile.scala 38:30]
  wire  _T_26 = io_rs1_addr != 5'h0; // @[regfile.scala 48:36]
  wire  _T_31 = io_rs2_addr != 5'h0; // @[regfile.scala 49:36]
  wire [31:0] regfile__T_27_data = mem_sparse_io_r_0_data;
  wire [31:0] regfile__T_32_data = mem_sparse_io_r_1_data;
  SparseMem mem_sparse (
    .metaReset(mem_sparse_metaReset),
    .clock(mem_sparse_clock),
    .io_w_0_addr(mem_sparse_io_w_0_addr),
    .io_w_0_en(mem_sparse_io_w_0_en),
    .io_w_0_data(mem_sparse_io_w_0_data),
    .io_r_0_addr(mem_sparse_io_r_0_addr),
    .io_r_0_data(mem_sparse_io_r_0_data),
    .io_r_1_addr(mem_sparse_io_r_1_addr),
    .io_r_1_data(mem_sparse_io_r_1_data)
  );
  assign mem_sparse_metaReset = metaReset;
  assign io_rs1_data = _T_26 ? regfile__T_27_data : 32'h0; // @[regfile.scala 48:16]
  assign io_rs2_data = _T_31 ? regfile__T_32_data : 32'h0; // @[regfile.scala 49:16]
  assign _GEN_0_0 = io_rs1_addr != 5'h0;
  assign _GEN_1_3 = io_rs2_addr != 5'h0;
  assign mem_sparse_clock = clock;
  assign mem_sparse_io_w_0_addr = io_waddr;
  assign mem_sparse_io_w_0_en = io_wen & _T_18;
  assign mem_sparse_io_w_0_data = io_wdata;
  assign mem_sparse_io_r_0_addr = io_rs1_addr;
  assign mem_sparse_io_r_1_addr = io_rs2_addr;
endmodule
module SparseMem(
  input         metaReset,
  input         clock,
  input  [4:0]  io_w_0_addr,
  input         io_w_0_en,
  input  [31:0] io_w_0_data,
  input  [4:0]  io_r_0_addr,
  output [31:0] io_r_0_data,
  input  [4:0]  io_r_1_addr,
  output [31:0] io_r_1_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:31];
  wire [31:0] mem__T_152_data;
  wire [4:0] mem__T_152_addr;
  wire [31:0] mem__T_274_data;
  wire [4:0] mem__T_274_addr;
  wire [31:0] mem__T_396_data;
  wire [4:0] mem__T_396_addr;
  wire [31:0] mem__T_528_data;
  wire [4:0] mem__T_528_addr;
  wire  mem__T_528_mask;
  wire  mem__T_528_en;
  wire [31:0] mem__T_656_data;
  wire [4:0] mem__T_656_addr;
  wire  mem__T_656_mask;
  wire  mem__T_656_en;
  reg [4:0] addresses_0_bits;
  reg [4:0] addresses_1_bits;
  reg [4:0] addresses_2_bits;
  reg [4:0] addresses_3_bits;
  reg [4:0] addresses_4_bits;
  reg [4:0] addresses_5_bits;
  reg [4:0] addresses_6_bits;
  reg [4:0] addresses_7_bits;
  reg [4:0] addresses_8_bits;
  reg [4:0] addresses_9_bits;
  reg [4:0] addresses_10_bits;
  reg [4:0] addresses_11_bits;
  reg [4:0] addresses_12_bits;
  reg [4:0] addresses_13_bits;
  reg [4:0] addresses_14_bits;
  reg [4:0] addresses_15_bits;
  reg [4:0] addresses_16_bits;
  reg [4:0] addresses_17_bits;
  reg [4:0] addresses_18_bits;
  reg [4:0] addresses_19_bits;
  reg [4:0] addresses_20_bits;
  reg [4:0] addresses_21_bits;
  reg [4:0] addresses_22_bits;
  reg [4:0] addresses_23_bits;
  reg [4:0] addresses_24_bits;
  reg [4:0] addresses_25_bits;
  reg [4:0] addresses_26_bits;
  reg [4:0] addresses_27_bits;
  reg [4:0] addresses_28_bits;
  reg [4:0] addresses_29_bits;
  reg [4:0] addresses_30_bits;
  reg [4:0] addresses_31_bits;
  wire  _T_33 = addresses_0_bits == io_r_0_addr;
  wire  _T_35 = addresses_1_bits == io_r_0_addr;
  wire  _T_37 = addresses_2_bits == io_r_0_addr;
  wire  _T_39 = addresses_3_bits == io_r_0_addr;
  wire  _T_41 = addresses_4_bits == io_r_0_addr;
  wire  _T_43 = addresses_5_bits == io_r_0_addr;
  wire  _T_45 = addresses_6_bits == io_r_0_addr;
  wire  _T_47 = addresses_7_bits == io_r_0_addr;
  wire  _T_49 = addresses_8_bits == io_r_0_addr;
  wire  _T_51 = addresses_9_bits == io_r_0_addr;
  wire  _T_53 = addresses_10_bits == io_r_0_addr;
  wire  _T_55 = addresses_11_bits == io_r_0_addr;
  wire  _T_57 = addresses_12_bits == io_r_0_addr;
  wire  _T_59 = addresses_13_bits == io_r_0_addr;
  wire  _T_61 = addresses_14_bits == io_r_0_addr;
  wire  _T_63 = addresses_15_bits == io_r_0_addr;
  wire  _T_65 = addresses_16_bits == io_r_0_addr;
  wire  _T_67 = addresses_17_bits == io_r_0_addr;
  wire  _T_69 = addresses_18_bits == io_r_0_addr;
  wire  _T_71 = addresses_19_bits == io_r_0_addr;
  wire  _T_73 = addresses_20_bits == io_r_0_addr;
  wire  _T_75 = addresses_21_bits == io_r_0_addr;
  wire  _T_77 = addresses_22_bits == io_r_0_addr;
  wire  _T_79 = addresses_23_bits == io_r_0_addr;
  wire  _T_81 = addresses_24_bits == io_r_0_addr;
  wire  _T_83 = addresses_25_bits == io_r_0_addr;
  wire  _T_85 = addresses_26_bits == io_r_0_addr;
  wire  _T_87 = addresses_27_bits == io_r_0_addr;
  wire  _T_89 = addresses_28_bits == io_r_0_addr;
  wire  _T_91 = addresses_29_bits == io_r_0_addr;
  wire  _T_93 = addresses_30_bits == io_r_0_addr;
  wire  _T_95 = addresses_31_bits == io_r_0_addr;
  wire [7:0] _T_104 = {_T_47,_T_45,_T_43,_T_41,_T_39,_T_37,_T_35,_T_33};
  wire [15:0] _T_112 = {_T_63,_T_61,_T_59,_T_57,_T_55,_T_53,_T_51,_T_49,_T_104};
  wire [7:0] _T_119 = {_T_79,_T_77,_T_75,_T_73,_T_71,_T_69,_T_67,_T_65};
  wire [31:0] _T_128 = {_T_95,_T_93,_T_91,_T_89,_T_87,_T_85,_T_83,_T_81,_T_119,_T_112};
  wire  _T_129 = _T_128 != 32'h0;
  wire  _T_132 = |_T_128[31:16];
  wire [15:0] _T_133 = _T_128[31:16] | _T_128[15:0];
  wire  _T_136 = |_T_133[15:8];
  wire [7:0] _T_137 = _T_133[15:8] | _T_133[7:0];
  wire  _T_140 = |_T_137[7:4];
  wire [3:0] _T_141 = _T_137[7:4] | _T_137[3:0];
  wire  _T_144 = |_T_141[3:2];
  wire [1:0] _T_145 = _T_141[3:2] | _T_141[1:0];
  wire [3:0] _T_149 = {_T_136,_T_140,_T_144,_T_145[1]};
  wire  _T_155 = addresses_0_bits == io_r_1_addr;
  wire  _T_157 = addresses_1_bits == io_r_1_addr;
  wire  _T_159 = addresses_2_bits == io_r_1_addr;
  wire  _T_161 = addresses_3_bits == io_r_1_addr;
  wire  _T_163 = addresses_4_bits == io_r_1_addr;
  wire  _T_165 = addresses_5_bits == io_r_1_addr;
  wire  _T_167 = addresses_6_bits == io_r_1_addr;
  wire  _T_169 = addresses_7_bits == io_r_1_addr;
  wire  _T_171 = addresses_8_bits == io_r_1_addr;
  wire  _T_173 = addresses_9_bits == io_r_1_addr;
  wire  _T_175 = addresses_10_bits == io_r_1_addr;
  wire  _T_177 = addresses_11_bits == io_r_1_addr;
  wire  _T_179 = addresses_12_bits == io_r_1_addr;
  wire  _T_181 = addresses_13_bits == io_r_1_addr;
  wire  _T_183 = addresses_14_bits == io_r_1_addr;
  wire  _T_185 = addresses_15_bits == io_r_1_addr;
  wire  _T_187 = addresses_16_bits == io_r_1_addr;
  wire  _T_189 = addresses_17_bits == io_r_1_addr;
  wire  _T_191 = addresses_18_bits == io_r_1_addr;
  wire  _T_193 = addresses_19_bits == io_r_1_addr;
  wire  _T_195 = addresses_20_bits == io_r_1_addr;
  wire  _T_197 = addresses_21_bits == io_r_1_addr;
  wire  _T_199 = addresses_22_bits == io_r_1_addr;
  wire  _T_201 = addresses_23_bits == io_r_1_addr;
  wire  _T_203 = addresses_24_bits == io_r_1_addr;
  wire  _T_205 = addresses_25_bits == io_r_1_addr;
  wire  _T_207 = addresses_26_bits == io_r_1_addr;
  wire  _T_209 = addresses_27_bits == io_r_1_addr;
  wire  _T_211 = addresses_28_bits == io_r_1_addr;
  wire  _T_213 = addresses_29_bits == io_r_1_addr;
  wire  _T_215 = addresses_30_bits == io_r_1_addr;
  wire  _T_217 = addresses_31_bits == io_r_1_addr;
  wire [7:0] _T_226 = {_T_169,_T_167,_T_165,_T_163,_T_161,_T_159,_T_157,_T_155};
  wire [15:0] _T_234 = {_T_185,_T_183,_T_181,_T_179,_T_177,_T_175,_T_173,_T_171,_T_226};
  wire [7:0] _T_241 = {_T_201,_T_199,_T_197,_T_195,_T_193,_T_191,_T_189,_T_187};
  wire [31:0] _T_250 = {_T_217,_T_215,_T_213,_T_211,_T_209,_T_207,_T_205,_T_203,_T_241,_T_234};
  wire  _T_251 = _T_250 != 32'h0;
  wire  _T_254 = |_T_250[31:16];
  wire [15:0] _T_255 = _T_250[31:16] | _T_250[15:0];
  wire  _T_258 = |_T_255[15:8];
  wire [7:0] _T_259 = _T_255[15:8] | _T_255[7:0];
  wire  _T_262 = |_T_259[7:4];
  wire [3:0] _T_263 = _T_259[7:4] | _T_259[3:0];
  wire  _T_266 = |_T_263[3:2];
  wire [1:0] _T_267 = _T_263[3:2] | _T_263[1:0];
  wire [3:0] _T_271 = {_T_258,_T_262,_T_266,_T_267[1]};
  wire  _T_277 = addresses_0_bits == 5'h0;
  wire  _T_279 = addresses_1_bits == 5'h0;
  wire  _T_281 = addresses_2_bits == 5'h0;
  wire  _T_283 = addresses_3_bits == 5'h0;
  wire  _T_285 = addresses_4_bits == 5'h0;
  wire  _T_287 = addresses_5_bits == 5'h0;
  wire  _T_289 = addresses_6_bits == 5'h0;
  wire  _T_291 = addresses_7_bits == 5'h0;
  wire  _T_293 = addresses_8_bits == 5'h0;
  wire  _T_295 = addresses_9_bits == 5'h0;
  wire  _T_297 = addresses_10_bits == 5'h0;
  wire  _T_299 = addresses_11_bits == 5'h0;
  wire  _T_301 = addresses_12_bits == 5'h0;
  wire  _T_303 = addresses_13_bits == 5'h0;
  wire  _T_305 = addresses_14_bits == 5'h0;
  wire  _T_307 = addresses_15_bits == 5'h0;
  wire  _T_309 = addresses_16_bits == 5'h0;
  wire  _T_311 = addresses_17_bits == 5'h0;
  wire  _T_313 = addresses_18_bits == 5'h0;
  wire  _T_315 = addresses_19_bits == 5'h0;
  wire  _T_317 = addresses_20_bits == 5'h0;
  wire  _T_319 = addresses_21_bits == 5'h0;
  wire  _T_321 = addresses_22_bits == 5'h0;
  wire  _T_323 = addresses_23_bits == 5'h0;
  wire  _T_325 = addresses_24_bits == 5'h0;
  wire  _T_327 = addresses_25_bits == 5'h0;
  wire  _T_329 = addresses_26_bits == 5'h0;
  wire  _T_331 = addresses_27_bits == 5'h0;
  wire  _T_333 = addresses_28_bits == 5'h0;
  wire  _T_335 = addresses_29_bits == 5'h0;
  wire  _T_337 = addresses_30_bits == 5'h0;
  wire  _T_339 = addresses_31_bits == 5'h0;
  wire [7:0] _T_348 = {_T_291,_T_289,_T_287,_T_285,_T_283,_T_281,_T_279,_T_277};
  wire [15:0] _T_356 = {_T_307,_T_305,_T_303,_T_301,_T_299,_T_297,_T_295,_T_293,_T_348};
  wire [7:0] _T_363 = {_T_323,_T_321,_T_319,_T_317,_T_315,_T_313,_T_311,_T_309};
  wire [31:0] _T_372 = {_T_339,_T_337,_T_335,_T_333,_T_331,_T_329,_T_327,_T_325,_T_363,_T_356};
  wire  _T_373 = _T_372 != 32'h0;
  wire  _T_376 = |_T_372[31:16];
  wire [15:0] _T_377 = _T_372[31:16] | _T_372[15:0];
  wire  _T_380 = |_T_377[15:8];
  wire [7:0] _T_381 = _T_377[15:8] | _T_377[7:0];
  wire  _T_384 = |_T_381[7:4];
  wire [3:0] _T_385 = _T_381[7:4] | _T_381[3:0];
  wire  _T_388 = |_T_385[3:2];
  wire [1:0] _T_389 = _T_385[3:2] | _T_385[1:0];
  wire [3:0] _T_393 = {_T_380,_T_384,_T_388,_T_389[1]};
  wire [4:0] _T_394 = {_T_376,_T_380,_T_384,_T_388,_T_389[1]};
  reg [5:0] nextAddr;
  wire [5:0] _T_400 = nextAddr + 6'h1;
  wire  _T_404 = addresses_0_bits == io_w_0_addr;
  wire  _T_406 = addresses_1_bits == io_w_0_addr;
  wire  _T_408 = addresses_2_bits == io_w_0_addr;
  wire  _T_410 = addresses_3_bits == io_w_0_addr;
  wire  _T_412 = addresses_4_bits == io_w_0_addr;
  wire  _T_414 = addresses_5_bits == io_w_0_addr;
  wire  _T_416 = addresses_6_bits == io_w_0_addr;
  wire  _T_418 = addresses_7_bits == io_w_0_addr;
  wire  _T_420 = addresses_8_bits == io_w_0_addr;
  wire  _T_422 = addresses_9_bits == io_w_0_addr;
  wire  _T_424 = addresses_10_bits == io_w_0_addr;
  wire  _T_426 = addresses_11_bits == io_w_0_addr;
  wire  _T_428 = addresses_12_bits == io_w_0_addr;
  wire  _T_430 = addresses_13_bits == io_w_0_addr;
  wire  _T_432 = addresses_14_bits == io_w_0_addr;
  wire  _T_434 = addresses_15_bits == io_w_0_addr;
  wire  _T_436 = addresses_16_bits == io_w_0_addr;
  wire  _T_438 = addresses_17_bits == io_w_0_addr;
  wire  _T_440 = addresses_18_bits == io_w_0_addr;
  wire  _T_442 = addresses_19_bits == io_w_0_addr;
  wire  _T_444 = addresses_20_bits == io_w_0_addr;
  wire  _T_446 = addresses_21_bits == io_w_0_addr;
  wire  _T_448 = addresses_22_bits == io_w_0_addr;
  wire  _T_450 = addresses_23_bits == io_w_0_addr;
  wire  _T_452 = addresses_24_bits == io_w_0_addr;
  wire  _T_454 = addresses_25_bits == io_w_0_addr;
  wire  _T_456 = addresses_26_bits == io_w_0_addr;
  wire  _T_458 = addresses_27_bits == io_w_0_addr;
  wire  _T_460 = addresses_28_bits == io_w_0_addr;
  wire  _T_462 = addresses_29_bits == io_w_0_addr;
  wire  _T_464 = addresses_30_bits == io_w_0_addr;
  wire  _T_466 = addresses_31_bits == io_w_0_addr;
  wire [7:0] _T_475 = {_T_418,_T_416,_T_414,_T_412,_T_410,_T_408,_T_406,_T_404};
  wire [15:0] _T_483 = {_T_434,_T_432,_T_430,_T_428,_T_426,_T_424,_T_422,_T_420,_T_475};
  wire [7:0] _T_490 = {_T_450,_T_448,_T_446,_T_444,_T_442,_T_440,_T_438,_T_436};
  wire [31:0] _T_499 = {_T_466,_T_464,_T_462,_T_460,_T_458,_T_456,_T_454,_T_452,_T_490,_T_483};
  wire  _T_500 = _T_499 != 32'h0;
  wire  _T_503 = |_T_499[31:16];
  wire [15:0] _T_504 = _T_499[31:16] | _T_499[15:0];
  wire  _T_507 = |_T_504[15:8];
  wire [7:0] _T_508 = _T_504[15:8] | _T_504[7:0];
  wire  _T_511 = |_T_508[7:4];
  wire [3:0] _T_512 = _T_508[7:4] | _T_508[3:0];
  wire  _T_515 = |_T_512[3:2];
  wire [1:0] _T_516 = _T_512[3:2] | _T_512[1:0];
  wire [4:0] _T_521 = {_T_503,_T_507,_T_511,_T_515,_T_516[1]};
  wire  _T_522 = ~_T_500;
  wire  _T_523 = io_w_0_en & _T_522;
  wire [5:0] _T_524 = _T_500 ? {{1'd0}, _T_521} : nextAddr;
  wire [5:0] nextAddrUpdate = _T_523 ? _T_400 : nextAddr;
  wire [5:0] _T_652 = _T_373 ? {{1'd0}, _T_394} : nextAddrUpdate;
  wire  _T_659 = nextAddrUpdate <= 6'h20;
  wire  _T_662 = ~_T_659;
  assign mem__T_152_addr = {_T_132,_T_149};
  assign mem__T_152_data = mem[mem__T_152_addr];
  assign mem__T_274_addr = {_T_254,_T_271};
  assign mem__T_274_data = mem[mem__T_274_addr];
  assign mem__T_396_addr = {_T_376,_T_393};
  assign mem__T_396_data = mem[mem__T_396_addr];
  assign mem__T_528_data = io_w_0_data;
  assign mem__T_528_addr = _T_524[4:0];
  assign mem__T_528_mask = 1'h1;
  assign mem__T_528_en = io_w_0_en;
  assign mem__T_656_data = 32'h0;
  assign mem__T_656_addr = _T_652[4:0];
  assign mem__T_656_mask = 1'h1;
  assign mem__T_656_en = 1'h0;
  assign io_r_0_data = _T_129 ? mem__T_152_data : 32'h0;
  assign io_r_1_data = _T_251 ? mem__T_274_data : 32'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  addresses_0_bits = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  addresses_1_bits = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  addresses_2_bits = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  addresses_3_bits = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  addresses_4_bits = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  addresses_5_bits = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  addresses_6_bits = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  addresses_7_bits = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  addresses_8_bits = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  addresses_9_bits = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  addresses_10_bits = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  addresses_11_bits = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  addresses_12_bits = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  addresses_13_bits = _RAND_14[4:0];
  _RAND_15 = {1{`RANDOM}};
  addresses_14_bits = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  addresses_15_bits = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  addresses_16_bits = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  addresses_17_bits = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  addresses_18_bits = _RAND_19[4:0];
  _RAND_20 = {1{`RANDOM}};
  addresses_19_bits = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  addresses_20_bits = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  addresses_21_bits = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  addresses_22_bits = _RAND_23[4:0];
  _RAND_24 = {1{`RANDOM}};
  addresses_23_bits = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  addresses_24_bits = _RAND_25[4:0];
  _RAND_26 = {1{`RANDOM}};
  addresses_25_bits = _RAND_26[4:0];
  _RAND_27 = {1{`RANDOM}};
  addresses_26_bits = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  addresses_27_bits = _RAND_28[4:0];
  _RAND_29 = {1{`RANDOM}};
  addresses_28_bits = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  addresses_29_bits = _RAND_30[4:0];
  _RAND_31 = {1{`RANDOM}};
  addresses_30_bits = _RAND_31[4:0];
  _RAND_32 = {1{`RANDOM}};
  addresses_31_bits = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  nextAddr = _RAND_33[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_528_en & mem__T_528_mask) begin
      mem[mem__T_528_addr] <= mem__T_528_data;
    end
    if(mem__T_656_en & mem__T_656_mask) begin
      mem[mem__T_656_addr] <= mem__T_656_data;
    end
    if (metaReset) begin
      addresses_0_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h0 == _T_524[4:0]) begin
        addresses_0_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_1_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h1 == _T_524[4:0]) begin
        addresses_1_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_2_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h2 == _T_524[4:0]) begin
        addresses_2_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_3_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h3 == _T_524[4:0]) begin
        addresses_3_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_4_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h4 == _T_524[4:0]) begin
        addresses_4_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_5_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h5 == _T_524[4:0]) begin
        addresses_5_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_6_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h6 == _T_524[4:0]) begin
        addresses_6_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_7_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h7 == _T_524[4:0]) begin
        addresses_7_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_8_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h8 == _T_524[4:0]) begin
        addresses_8_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_9_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h9 == _T_524[4:0]) begin
        addresses_9_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_10_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'ha == _T_524[4:0]) begin
        addresses_10_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_11_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'hb == _T_524[4:0]) begin
        addresses_11_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_12_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'hc == _T_524[4:0]) begin
        addresses_12_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_13_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'hd == _T_524[4:0]) begin
        addresses_13_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_14_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'he == _T_524[4:0]) begin
        addresses_14_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_15_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'hf == _T_524[4:0]) begin
        addresses_15_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_16_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h10 == _T_524[4:0]) begin
        addresses_16_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_17_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h11 == _T_524[4:0]) begin
        addresses_17_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_18_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h12 == _T_524[4:0]) begin
        addresses_18_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_19_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h13 == _T_524[4:0]) begin
        addresses_19_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_20_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h14 == _T_524[4:0]) begin
        addresses_20_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_21_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h15 == _T_524[4:0]) begin
        addresses_21_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_22_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h16 == _T_524[4:0]) begin
        addresses_22_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_23_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h17 == _T_524[4:0]) begin
        addresses_23_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_24_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h18 == _T_524[4:0]) begin
        addresses_24_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_25_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h19 == _T_524[4:0]) begin
        addresses_25_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_26_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h1a == _T_524[4:0]) begin
        addresses_26_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_27_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h1b == _T_524[4:0]) begin
        addresses_27_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_28_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h1c == _T_524[4:0]) begin
        addresses_28_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_29_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h1d == _T_524[4:0]) begin
        addresses_29_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_30_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h1e == _T_524[4:0]) begin
        addresses_30_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      addresses_31_bits <= 5'h0;
    end else if (io_w_0_en) begin
      if (5'h1f == _T_524[4:0]) begin
        addresses_31_bits <= io_w_0_addr;
      end
    end
    if (metaReset) begin
      nextAddr <= 6'h0;
    end else if (_T_523) begin
      nextAddr <= _T_400;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CSRFile(
  input         metaReset,
  input         clock,
  input         reset,
  input  [2:0]  io_rw_cmd,
  output [31:0] io_rw_rdata,
  input  [31:0] io_rw_wdata,
  output        io_eret,
  input  [11:0] io_decode_csr,
  output        io_status_debug,
  output [1:0]  io_status_prv,
  output        io_status_sd,
  output [7:0]  io_status_zero1,
  output        io_status_tsr,
  output        io_status_tw,
  output        io_status_tvm,
  output        io_status_mxr,
  output        io_status_sum,
  output        io_status_mprv,
  output [1:0]  io_status_xs,
  output [1:0]  io_status_fs,
  output [1:0]  io_status_mpp,
  output [1:0]  io_status_hpp,
  output        io_status_spp,
  output        io_status_mpie,
  output        io_status_hpie,
  output        io_status_spie,
  output        io_status_upie,
  output        io_status_mie,
  output        io_status_hie,
  output        io_status_sie,
  output        io_status_uie,
  output [31:0] io_evec,
  input         io_exception,
  input         io_retire,
  input  [31:0] io_pc,
  output        _GEN_451_0,
  output        _GEN_331_0,
  output        _GEN_337_0,
  output        _GEN_415_0,
  output        _GEN_436_0,
  output        _GEN_352_0,
  output        _GEN_430_0,
  output        _GEN_151_0,
  output        _GEN_310_0,
  output        _GEN_409_0,
  output        _GEN_253_0,
  output        _GEN_316_0,
  output        _GEN_244_0,
  output        _GEN_238_0,
  output        _GEN_325_0,
  output        _GEN_433_0,
  output        _GEN_313_0,
  output        _GEN_11_0,
  output        _GEN_304_0,
  output        _GEN_294_0,
  output        _GEN_303_0,
  output        _GEN_402_0,
  output        _GEN_412_0,
  output        _GEN_424_0,
  output        _GEN_319_0,
  output        _GEN_288_0,
  output        _GEN_418_0,
  output        _GEN_387_0,
  output        _GEN_462_0,
  output        _GEN_375_0,
  output        _GEN_390_0,
  output        _GEN_307_0,
  output        _GEN_297_0,
  output        _GEN_406_0,
  output        _GEN_270_0,
  output        _GEN_369_0,
  output        _GEN_396_0,
  output        _GEN_276_0,
  output        _GEN_291_0,
  output        _GEN_258_0,
  output        _GEN_372_0,
  output        _GEN_252_1,
  output        _GEN_285_0,
  output        _GEN_384_0,
  output        _GEN_378_0,
  output        _GEN_393_0,
  output        _GEN_273_0,
  output        _GEN_456_0,
  output        _GEN_351_1,
  output        _GEN_450_0,
  output        _GEN_357_0,
  output        _GEN_279_0,
  output        _GEN_399_0,
  output        _GEN_264_0,
  output        _GEN_300_0,
  output        _GEN_432_0,
  output        _GEN_381_0,
  output        _GEN_339_1,
  output        _GEN_261_0,
  output        _GEN_360_0,
  output        _GEN_246_1,
  output        _GEN_438_0,
  output        _GEN_282_0,
  output        _GEN_345_1,
  output        _GEN_240_1,
  output        _GEN_444_0,
  output        _GEN_267_1,
  output        _GEN_459_0,
  output        _GEN_453_0,
  output        _GEN_366_0,
  output        _GEN_7_0,
  output        _GEN_324_1,
  output        _GEN_333_1,
  output        _GEN_342_0,
  output        _GEN_405_0,
  output        _GEN_420_1,
  output        _GEN_306_0,
  output        _GEN_3_0,
  output        _GEN_426_0,
  output        _GEN_441_0,
  output        _GEN_348_0,
  output        _GEN_255_0,
  output        _GEN_146_0,
  output        _GEN_363_0,
  output        _GEN_321_1,
  output        _GEN_327_1,
  output        _GEN_354_0,
  output        _GEN_234_1,
  output        _GEN_249_1,
  output        _GEN_243_0,
  output        _GEN_447_0,
  output        _GEN_330_1,
  output        _GEN_429_0,
  output        _GEN_293_1,
  output        _GEN_414_1,
  output        _GEN_309_0,
  output        _GEN_299_1,
  output        _GEN_336_0,
  output        _GEN_408_0,
  output        _GEN_150_0,
  output        _GEN_435_0,
  output        _GEN_392_1,
  output        _GEN_398_1,
  output        _GEN_423_1,
  output        _GEN_237_0,
  output        _GEN_315_1,
  output        _GEN_302_1,
  output        _GEN_380_1,
  output        _GEN_318_1,
  output        _GEN_287_1,
  output        _GEN_386_1,
  output        _GEN_281_1,
  output        _GEN_312_1,
  output        _GEN_417_1,
  output        _GEN_411_1,
  output        _GEN_401_1,
  output        _GEN_374_1,
  output        _GEN_368_1,
  output        _GEN_383_1,
  output        _GEN_263_1,
  output        _GEN_446_0,
  output        _GEN_290_1,
  output        _GEN_389_1,
  output        _GEN_254_1,
  output        _GEN_461_0,
  output        _GEN_362_1,
  output        _GEN_296_1,
  output        _GEN_395_1,
  output        _GEN_275_1,
  output        _GEN_269_1,
  output        _GEN_278_1,
  output        _GEN_251_1,
  output        _GEN_455_0,
  output        _GEN_377_1,
  output        _GEN_272_1,
  output        _GEN_335_1,
  output        _GEN_434_0,
  output        _GEN_257_1,
  output        _GEN_443_0,
  output        _GEN_356_1,
  output        _GEN_350_1,
  output        _GEN_428_0,
  output        _GEN_449_0,
  output        _GEN_236_1,
  output        _GEN_371_1,
  output        _GEN_284_1,
  output        _GEN_416_1,
  output        _GEN_260_1,
  output        _GEN_338_1,
  output        _GEN_344_1,
  output        _GEN_239_1,
  output        _GEN_353_1,
  output        _GEN_266_1,
  output        _GEN_452_0,
  output        _GEN_365_1,
  output        _GEN_6_0,
  output        _GEN_410_1,
  output        _GEN_152_1,
  output        _GEN_437_0,
  output        _GEN_332_1,
  output        _GEN_245_1,
  output        _GEN_359_1,
  output        _GEN_431_0,
  output        _GEN_458_0,
  output        _GEN_317_1,
  output        _GEN_326_1,
  output        _GEN_341_1,
  output        _GEN_394_1,
  output        _GEN_248_1,
  output        _GEN_347_1,
  output        _GEN_425_1,
  output        _GEN_305_1,
  output        _GEN_419_1,
  output        _GEN_320_1,
  output        _GEN_413_1,
  output        _GEN_440_0,
  output        _GEN_295_1,
  output        _GEN_404_1,
  output        _GEN_403_1,
  output        _GEN_242_1,
  output        _GEN_15_1,
  output        _GEN_308_1,
  output        _GEN_149_1,
  output        _GEN_329_1,
  output        _GEN_292_1,
  output        _GEN_298_1,
  output        _GEN_391_1,
  output        _GEN_314_1,
  output        _GEN_323_1,
  output        _GEN_376_1,
  output        _GEN_422_1,
  output        _GEN_277_1,
  output        _GEN_407_1,
  output        _GEN_397_1,
  output        _GEN_379_1,
  output        _GEN_373_1,
  output        _GEN_364_1,
  output        _GEN_259_1,
  output        _GEN_265_1,
  output        _GEN_301_1,
  output        _GEN_286_1,
  output        _GEN_400_1,
  output        _GEN_358_1,
  output        _GEN_385_1,
  output        _GEN_457_0,
  output        _GEN_311_1,
  output        _GEN_280_1,
  output        _GEN_367_1,
  output        _GEN_247_1,
  output        _GEN_274_1,
  output        _GEN_460_0,
  output        _GEN_283_1,
  output        _GEN_388_1,
  output        _GEN_382_1,
  output        _GEN_268_1,
  output        _GEN_346_1,
  output        _GEN_340_1,
  output        _GEN_439_0,
  output        _GEN_262_1,
  output        _GEN_361_1,
  output        _GEN_241_1,
  output        _GEN_445_0,
  output        _GEN_289_1,
  output        _GEN_421_1,
  output        _GEN_427_0,
  output        _GEN_454_0,
  output        _GEN_256_1,
  output        _GEN_5_2,
  output        _GEN_271_1,
  output        _GEN_322_1,
  output        _GEN_334_1,
  output        _GEN_235_1,
  output        _GEN_349_1,
  output        _GEN_147_2,
  output        _GEN_448_0,
  output        _GEN_442_0,
  output        _GEN_343_1,
  output        _GEN_355_1,
  output        _GEN_370_1,
  output        _GEN_250_1,
  output        _GEN_463_0,
  output        _GEN_328_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
`endif // RANDOMIZE_REG_INIT
  reg  reg_mstatus_mpie; // @[csr.scala 163:24]
  reg  reg_mstatus_mie; // @[csr.scala 163:24]
  reg [31:0] reg_mepc; // @[csr.scala 164:21]
  reg [31:0] reg_mcause; // @[csr.scala 165:23]
  reg [31:0] reg_mtval; // @[csr.scala 166:22]
  reg [31:0] reg_mscratch; // @[csr.scala 167:25]
  reg [31:0] reg_medeleg; // @[csr.scala 169:24]
  reg  reg_mip_mtip; // @[csr.scala 171:20]
  reg  reg_mip_msip; // @[csr.scala 171:20]
  reg  reg_mie_mtip; // @[csr.scala 172:20]
  reg  reg_mie_msip; // @[csr.scala 172:20]
  reg [5:0] _T_176; // @[util.scala 114:37]
  wire [6:0] _T_177 = _T_176 + 6'h1; // @[util.scala 115:33]
  reg [57:0] _T_180; // @[util.scala 119:27]
  wire [57:0] _T_184 = _T_180 + 58'h1; // @[util.scala 120:43]
  wire [63:0] _T_185 = {_T_180,_T_176}; // @[Cat.scala 30:58]
  reg [5:0] _T_188; // @[util.scala 114:37]
  wire [5:0] _GEN_153 = {{5'd0}, io_retire}; // @[util.scala 115:33]
  wire [6:0] _T_189 = _T_188 + _GEN_153; // @[util.scala 115:33]
  reg [57:0] _T_192; // @[util.scala 119:27]
  wire [57:0] _T_196 = _T_192 + 58'h1; // @[util.scala 120:43]
  wire [63:0] _T_197 = {_T_192,_T_188}; // @[Cat.scala 30:58]
  reg [39:0] _T_200; // @[util.scala 114:75]
  wire [40:0] _T_201 = {{1'd0}, _T_200}; // @[util.scala 115:33]
  reg [39:0] _T_203; // @[util.scala 114:75]
  wire [40:0] _T_204 = {{1'd0}, _T_203}; // @[util.scala 115:33]
  reg [39:0] _T_206; // @[util.scala 114:75]
  wire [40:0] _T_207 = {{1'd0}, _T_206}; // @[util.scala 115:33]
  reg [39:0] _T_209; // @[util.scala 114:75]
  wire [40:0] _T_210 = {{1'd0}, _T_209}; // @[util.scala 115:33]
  reg [39:0] _T_212; // @[util.scala 114:75]
  wire [40:0] _T_213 = {{1'd0}, _T_212}; // @[util.scala 115:33]
  reg [39:0] _T_215; // @[util.scala 114:75]
  wire [40:0] _T_216 = {{1'd0}, _T_215}; // @[util.scala 115:33]
  reg [39:0] _T_218; // @[util.scala 114:75]
  wire [40:0] _T_219 = {{1'd0}, _T_218}; // @[util.scala 115:33]
  reg [39:0] _T_221; // @[util.scala 114:75]
  wire [40:0] _T_222 = {{1'd0}, _T_221}; // @[util.scala 115:33]
  reg [39:0] _T_224; // @[util.scala 114:75]
  wire [40:0] _T_225 = {{1'd0}, _T_224}; // @[util.scala 115:33]
  reg [39:0] _T_227; // @[util.scala 114:75]
  wire [40:0] _T_228 = {{1'd0}, _T_227}; // @[util.scala 115:33]
  reg [39:0] _T_230; // @[util.scala 114:75]
  wire [40:0] _T_231 = {{1'd0}, _T_230}; // @[util.scala 115:33]
  reg [39:0] _T_233; // @[util.scala 114:75]
  wire [40:0] _T_234 = {{1'd0}, _T_233}; // @[util.scala 115:33]
  reg [39:0] _T_236; // @[util.scala 114:75]
  wire [40:0] _T_237 = {{1'd0}, _T_236}; // @[util.scala 115:33]
  reg [39:0] _T_239; // @[util.scala 114:75]
  wire [40:0] _T_240 = {{1'd0}, _T_239}; // @[util.scala 115:33]
  reg [39:0] _T_242; // @[util.scala 114:75]
  wire [40:0] _T_243 = {{1'd0}, _T_242}; // @[util.scala 115:33]
  reg [39:0] _T_245; // @[util.scala 114:75]
  wire [40:0] _T_246 = {{1'd0}, _T_245}; // @[util.scala 115:33]
  reg [39:0] _T_248; // @[util.scala 114:75]
  wire [40:0] _T_249 = {{1'd0}, _T_248}; // @[util.scala 115:33]
  reg [39:0] _T_251; // @[util.scala 114:75]
  wire [40:0] _T_252 = {{1'd0}, _T_251}; // @[util.scala 115:33]
  reg [39:0] _T_254; // @[util.scala 114:75]
  wire [40:0] _T_255 = {{1'd0}, _T_254}; // @[util.scala 115:33]
  reg [39:0] _T_257; // @[util.scala 114:75]
  wire [40:0] _T_258 = {{1'd0}, _T_257}; // @[util.scala 115:33]
  reg [39:0] _T_260; // @[util.scala 114:75]
  wire [40:0] _T_261 = {{1'd0}, _T_260}; // @[util.scala 115:33]
  reg [39:0] _T_263; // @[util.scala 114:75]
  wire [40:0] _T_264 = {{1'd0}, _T_263}; // @[util.scala 115:33]
  reg [39:0] _T_266; // @[util.scala 114:75]
  wire [40:0] _T_267 = {{1'd0}, _T_266}; // @[util.scala 115:33]
  reg [39:0] _T_269; // @[util.scala 114:75]
  wire [40:0] _T_270 = {{1'd0}, _T_269}; // @[util.scala 115:33]
  reg [39:0] _T_272; // @[util.scala 114:75]
  wire [40:0] _T_273 = {{1'd0}, _T_272}; // @[util.scala 115:33]
  reg [39:0] _T_275; // @[util.scala 114:75]
  wire [40:0] _T_276 = {{1'd0}, _T_275}; // @[util.scala 115:33]
  reg [39:0] _T_278; // @[util.scala 114:75]
  wire [40:0] _T_279 = {{1'd0}, _T_278}; // @[util.scala 115:33]
  reg [39:0] _T_281; // @[util.scala 114:75]
  wire [40:0] _T_282 = {{1'd0}, _T_281}; // @[util.scala 115:33]
  reg [39:0] _T_284; // @[util.scala 114:75]
  wire [40:0] _T_285 = {{1'd0}, _T_284}; // @[util.scala 115:33]
  reg [39:0] _T_287; // @[util.scala 114:75]
  wire [40:0] _T_288 = {{1'd0}, _T_287}; // @[util.scala 115:33]
  reg [39:0] _T_290; // @[util.scala 114:75]
  wire [40:0] _T_291 = {{1'd0}, _T_290}; // @[util.scala 115:33]
  reg [39:0] _T_293; // @[util.scala 114:75]
  wire [40:0] _T_294 = {{1'd0}, _T_293}; // @[util.scala 115:33]
  reg [31:0] reg_dpc; // @[csr.scala 188:20]
  reg [31:0] reg_dscratch; // @[csr.scala 189:25]
  reg  reg_dcsr_ebreakm; // @[csr.scala 194:21]
  reg  reg_dcsr_step; // @[csr.scala 194:21]
  wire  system_insn = io_rw_cmd == 3'h4; // @[csr.scala 196:31]
  wire  _T_410 = io_rw_cmd != 3'h0; // @[csr.scala 197:27]
  wire  _T_412 = ~system_insn; // @[csr.scala 197:39]
  wire  cpu_ren = _T_410 & _T_412; // @[csr.scala 197:36]
  wire [4:0] _T_416 = {io_status_upie,io_status_mie,io_status_hie,io_status_sie,io_status_uie};
  wire [12:0] _T_422 = {io_status_mpp,io_status_hpp,io_status_spp,io_status_mpie,io_status_hpie,io_status_spie,_T_416};
  wire [7:0] _T_427 = {io_status_tvm,io_status_mxr,io_status_sum,io_status_mprv,io_status_xs,io_status_fs};
  wire [34:0] read_mstatus = {io_status_debug,io_status_prv,io_status_sd,io_status_zero1,io_status_tsr,io_status_tw,_T_427,_T_422};
  wire [15:0] _T_454 = {8'h0,reg_mip_mtip,1'h0,2'h0,reg_mip_msip,1'h0,2'h0};
  wire [15:0] _T_469 = {8'h0,reg_mie_mtip,1'h0,2'h0,reg_mie_msip,1'h0,2'h0};
  wire [31:0] _T_483 = {4'h4,12'h0,reg_dcsr_ebreakm,4'h0,6'h0,2'h0,reg_dcsr_step,2'h3}; // @[csr.scala 222:27]
  wire  _T_487 = io_decode_csr == 12'hb00; // @[csr.scala 259:76]
  wire  _T_489 = io_decode_csr == 12'hb02; // @[csr.scala 259:76]
  wire  _T_491 = io_decode_csr == 12'hf13; // @[csr.scala 259:76]
  wire  _T_497 = io_decode_csr == 12'h301; // @[csr.scala 259:76]
  wire  _T_499 = io_decode_csr == 12'h300; // @[csr.scala 259:76]
  wire  _T_501 = io_decode_csr == 12'h305; // @[csr.scala 259:76]
  wire  _T_503 = io_decode_csr == 12'h344; // @[csr.scala 259:76]
  wire  _T_505 = io_decode_csr == 12'h304; // @[csr.scala 259:76]
  wire  _T_507 = io_decode_csr == 12'h340; // @[csr.scala 259:76]
  wire  _T_509 = io_decode_csr == 12'h341; // @[csr.scala 259:76]
  wire  _T_511 = io_decode_csr == 12'h343; // @[csr.scala 259:76]
  wire  _T_513 = io_decode_csr == 12'h342; // @[csr.scala 259:76]
  wire  _T_517 = io_decode_csr == 12'h7b0; // @[csr.scala 259:76]
  wire  _T_519 = io_decode_csr == 12'h7b1; // @[csr.scala 259:76]
  wire  _T_521 = io_decode_csr == 12'h7b2; // @[csr.scala 259:76]
  wire  _T_523 = io_decode_csr == 12'h302; // @[csr.scala 259:76]
  wire  _T_525 = io_decode_csr == 12'hb03; // @[csr.scala 259:76]
  wire  _T_527 = io_decode_csr == 12'hb83; // @[csr.scala 259:76]
  wire  _T_529 = io_decode_csr == 12'hb04; // @[csr.scala 259:76]
  wire  _T_531 = io_decode_csr == 12'hb84; // @[csr.scala 259:76]
  wire  _T_533 = io_decode_csr == 12'hb05; // @[csr.scala 259:76]
  wire  _T_535 = io_decode_csr == 12'hb85; // @[csr.scala 259:76]
  wire  _T_537 = io_decode_csr == 12'hb06; // @[csr.scala 259:76]
  wire  _T_539 = io_decode_csr == 12'hb86; // @[csr.scala 259:76]
  wire  _T_541 = io_decode_csr == 12'hb07; // @[csr.scala 259:76]
  wire  _T_543 = io_decode_csr == 12'hb87; // @[csr.scala 259:76]
  wire  _T_545 = io_decode_csr == 12'hb08; // @[csr.scala 259:76]
  wire  _T_547 = io_decode_csr == 12'hb88; // @[csr.scala 259:76]
  wire  _T_549 = io_decode_csr == 12'hb09; // @[csr.scala 259:76]
  wire  _T_551 = io_decode_csr == 12'hb89; // @[csr.scala 259:76]
  wire  _T_553 = io_decode_csr == 12'hb0a; // @[csr.scala 259:76]
  wire  _T_555 = io_decode_csr == 12'hb8a; // @[csr.scala 259:76]
  wire  _T_557 = io_decode_csr == 12'hb0b; // @[csr.scala 259:76]
  wire  _T_559 = io_decode_csr == 12'hb8b; // @[csr.scala 259:76]
  wire  _T_561 = io_decode_csr == 12'hb0c; // @[csr.scala 259:76]
  wire  _T_563 = io_decode_csr == 12'hb8c; // @[csr.scala 259:76]
  wire  _T_565 = io_decode_csr == 12'hb0d; // @[csr.scala 259:76]
  wire  _T_567 = io_decode_csr == 12'hb8d; // @[csr.scala 259:76]
  wire  _T_569 = io_decode_csr == 12'hb0e; // @[csr.scala 259:76]
  wire  _T_571 = io_decode_csr == 12'hb8e; // @[csr.scala 259:76]
  wire  _T_573 = io_decode_csr == 12'hb0f; // @[csr.scala 259:76]
  wire  _T_575 = io_decode_csr == 12'hb8f; // @[csr.scala 259:76]
  wire  _T_577 = io_decode_csr == 12'hb10; // @[csr.scala 259:76]
  wire  _T_579 = io_decode_csr == 12'hb90; // @[csr.scala 259:76]
  wire  _T_581 = io_decode_csr == 12'hb11; // @[csr.scala 259:76]
  wire  _T_583 = io_decode_csr == 12'hb91; // @[csr.scala 259:76]
  wire  _T_585 = io_decode_csr == 12'hb12; // @[csr.scala 259:76]
  wire  _T_587 = io_decode_csr == 12'hb92; // @[csr.scala 259:76]
  wire  _T_589 = io_decode_csr == 12'hb13; // @[csr.scala 259:76]
  wire  _T_591 = io_decode_csr == 12'hb93; // @[csr.scala 259:76]
  wire  _T_593 = io_decode_csr == 12'hb14; // @[csr.scala 259:76]
  wire  _T_595 = io_decode_csr == 12'hb94; // @[csr.scala 259:76]
  wire  _T_597 = io_decode_csr == 12'hb15; // @[csr.scala 259:76]
  wire  _T_599 = io_decode_csr == 12'hb95; // @[csr.scala 259:76]
  wire  _T_601 = io_decode_csr == 12'hb16; // @[csr.scala 259:76]
  wire  _T_603 = io_decode_csr == 12'hb96; // @[csr.scala 259:76]
  wire  _T_605 = io_decode_csr == 12'hb17; // @[csr.scala 259:76]
  wire  _T_607 = io_decode_csr == 12'hb97; // @[csr.scala 259:76]
  wire  _T_609 = io_decode_csr == 12'hb18; // @[csr.scala 259:76]
  wire  _T_611 = io_decode_csr == 12'hb98; // @[csr.scala 259:76]
  wire  _T_613 = io_decode_csr == 12'hb19; // @[csr.scala 259:76]
  wire  _T_615 = io_decode_csr == 12'hb99; // @[csr.scala 259:76]
  wire  _T_617 = io_decode_csr == 12'hb1a; // @[csr.scala 259:76]
  wire  _T_619 = io_decode_csr == 12'hb9a; // @[csr.scala 259:76]
  wire  _T_621 = io_decode_csr == 12'hb1b; // @[csr.scala 259:76]
  wire  _T_623 = io_decode_csr == 12'hb9b; // @[csr.scala 259:76]
  wire  _T_625 = io_decode_csr == 12'hb1c; // @[csr.scala 259:76]
  wire  _T_627 = io_decode_csr == 12'hb9c; // @[csr.scala 259:76]
  wire  _T_629 = io_decode_csr == 12'hb1d; // @[csr.scala 259:76]
  wire  _T_631 = io_decode_csr == 12'hb9d; // @[csr.scala 259:76]
  wire  _T_633 = io_decode_csr == 12'hb1e; // @[csr.scala 259:76]
  wire  _T_635 = io_decode_csr == 12'hb9e; // @[csr.scala 259:76]
  wire  _T_637 = io_decode_csr == 12'hb1f; // @[csr.scala 259:76]
  wire  _T_639 = io_decode_csr == 12'hb9f; // @[csr.scala 259:76]
  wire  _T_641 = io_decode_csr == 12'hb20; // @[csr.scala 259:76]
  wire  _T_643 = io_decode_csr == 12'hba0; // @[csr.scala 259:76]
  wire  _T_645 = io_decode_csr == 12'hb21; // @[csr.scala 259:76]
  wire  _T_647 = io_decode_csr == 12'hba1; // @[csr.scala 259:76]
  wire  _T_649 = io_decode_csr == 12'hb22; // @[csr.scala 259:76]
  wire  _T_651 = io_decode_csr == 12'hba2; // @[csr.scala 259:76]
  wire  _T_653 = io_decode_csr == 12'hb80; // @[csr.scala 259:76]
  wire  _T_655 = io_decode_csr == 12'hb82; // @[csr.scala 259:76]
  wire [1:0] _T_658 = ~io_decode_csr[11:10]; // @[csr.scala 262:40]
  wire  read_only = _T_658 == 2'h0; // @[csr.scala 262:40]
  wire  _T_660 = io_rw_cmd != 3'h5; // @[csr.scala 263:38]
  wire  cpu_wen = cpu_ren & _T_660; // @[csr.scala 263:25]
  wire  _T_663 = ~read_only; // @[csr.scala 264:24]
  wire  wen = cpu_wen & _T_663; // @[csr.scala 264:21]
  wire  _T_664 = io_rw_cmd == 3'h2; // @[util.scala 25:47]
  wire  _T_665 = io_rw_cmd == 3'h3; // @[util.scala 25:47]
  wire  _T_666 = _T_664 | _T_665; // @[util.scala 25:62]
  wire [31:0] _T_668 = _T_666 ? io_rw_rdata : 32'h0; // @[csr.scala 390:9]
  wire [31:0] _T_669 = _T_668 | io_rw_wdata; // @[csr.scala 390:53]
  wire [31:0] _T_672 = _T_665 ? io_rw_wdata : 32'h0; // @[csr.scala 390:68]
  wire [31:0] _T_673 = ~_T_672; // @[csr.scala 390:64]
  wire [31:0] wdata = _T_669 & _T_673; // @[csr.scala 390:62]
  wire [7:0] opcode = 8'h1 << io_decode_csr[2:0]; // @[csr.scala 267:20]
  wire  insn_call = system_insn & opcode[0]; // @[csr.scala 268:31]
  wire  insn_break = system_insn & opcode[1]; // @[csr.scala 269:32]
  wire  insn_ret = system_insn & opcode[2]; // @[csr.scala 270:30]
  wire  _T_962 = insn_call | insn_break; // @[csr.scala 282:24]
  wire [31:0] _GEN_4 = io_exception ? io_pc : reg_mepc; // @[csr.scala 285:23]
  wire [1:0] _T_966 = insn_ret + io_exception; // @[Bitwise.scala 48:55]
  wire  _T_968 = _T_966 <= 2'h1; // @[csr.scala 291:52]
  wire  _T_970 = _T_968 | reset; // @[csr.scala 291:9]
  wire  _T_976 = insn_ret & io_decode_csr[10]; // @[csr.scala 298:17]
  wire [31:0] _GEN_8 = _T_976 ? reg_dpc : 32'h80000004; // @[csr.scala 298:38]
  wire  _T_980 = ~io_decode_csr[10]; // @[csr.scala 305:21]
  wire  _T_981 = insn_ret & _T_980; // @[csr.scala 305:18]
  wire  _GEN_10 = _T_981 | reg_mstatus_mpie; // @[csr.scala 305:41]
  wire [31:0] _GEN_12 = _T_981 ? reg_mepc : _GEN_8; // @[csr.scala 305:41]
  wire [31:0] _GEN_13 = insn_call ? 32'h80000004 : _GEN_12; // @[csr.scala 313:18]
  wire [63:0] _T_991 = _T_487 ? _T_185 : 64'h0; // @[Mux.scala 19:72]
  wire [63:0] _T_993 = _T_489 ? _T_197 : 64'h0; // @[Mux.scala 19:72]
  wire [15:0] _T_995 = _T_491 ? 16'h8000 : 16'h0; // @[Mux.scala 19:72]
  wire [8:0] _T_1001 = _T_497 ? 9'h100 : 9'h0; // @[Mux.scala 19:72]
  wire [34:0] _T_1003 = _T_499 ? read_mstatus : 35'h0; // @[Mux.scala 19:72]
  wire [8:0] _T_1005 = _T_501 ? 9'h100 : 9'h0; // @[Mux.scala 19:72]
  wire [15:0] _T_1007 = _T_503 ? _T_454 : 16'h0; // @[Mux.scala 19:72]
  wire [15:0] _T_1009 = _T_505 ? _T_469 : 16'h0; // @[Mux.scala 19:72]
  wire [31:0] _T_1011 = _T_507 ? reg_mscratch : 32'h0; // @[Mux.scala 19:72]
  wire [31:0] _T_1013 = _T_509 ? reg_mepc : 32'h0; // @[Mux.scala 19:72]
  wire [31:0] _T_1015 = _T_511 ? reg_mtval : 32'h0; // @[Mux.scala 19:72]
  wire [31:0] _T_1017 = _T_513 ? reg_mcause : 32'h0; // @[Mux.scala 19:72]
  wire [31:0] _T_1021 = _T_517 ? _T_483 : 32'h0; // @[Mux.scala 19:72]
  wire [31:0] _T_1023 = _T_519 ? reg_dpc : 32'h0; // @[Mux.scala 19:72]
  wire [31:0] _T_1025 = _T_521 ? reg_dscratch : 32'h0; // @[Mux.scala 19:72]
  wire [31:0] _T_1027 = _T_523 ? reg_medeleg : 32'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1029 = _T_525 ? _T_200 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1031 = _T_527 ? _T_200 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1033 = _T_529 ? _T_203 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1035 = _T_531 ? _T_203 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1037 = _T_533 ? _T_206 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1039 = _T_535 ? _T_206 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1041 = _T_537 ? _T_209 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1043 = _T_539 ? _T_209 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1045 = _T_541 ? _T_212 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1047 = _T_543 ? _T_212 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1049 = _T_545 ? _T_215 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1051 = _T_547 ? _T_215 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1053 = _T_549 ? _T_218 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1055 = _T_551 ? _T_218 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1057 = _T_553 ? _T_221 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1059 = _T_555 ? _T_221 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1061 = _T_557 ? _T_224 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1063 = _T_559 ? _T_224 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1065 = _T_561 ? _T_227 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1067 = _T_563 ? _T_227 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1069 = _T_565 ? _T_230 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1071 = _T_567 ? _T_230 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1073 = _T_569 ? _T_233 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1075 = _T_571 ? _T_233 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1077 = _T_573 ? _T_236 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1079 = _T_575 ? _T_236 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1081 = _T_577 ? _T_239 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1083 = _T_579 ? _T_239 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1085 = _T_581 ? _T_242 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1087 = _T_583 ? _T_242 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1089 = _T_585 ? _T_245 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1091 = _T_587 ? _T_245 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1093 = _T_589 ? _T_248 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1095 = _T_591 ? _T_248 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1097 = _T_593 ? _T_251 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1099 = _T_595 ? _T_251 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1101 = _T_597 ? _T_254 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1103 = _T_599 ? _T_254 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1105 = _T_601 ? _T_257 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1107 = _T_603 ? _T_257 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1109 = _T_605 ? _T_260 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1111 = _T_607 ? _T_260 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1113 = _T_609 ? _T_263 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1115 = _T_611 ? _T_263 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1117 = _T_613 ? _T_266 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1119 = _T_615 ? _T_266 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1121 = _T_617 ? _T_269 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1123 = _T_619 ? _T_269 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1125 = _T_621 ? _T_272 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1127 = _T_623 ? _T_272 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1129 = _T_625 ? _T_275 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1131 = _T_627 ? _T_275 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1133 = _T_629 ? _T_278 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1135 = _T_631 ? _T_278 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1137 = _T_633 ? _T_281 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1139 = _T_635 ? _T_281 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1141 = _T_637 ? _T_284 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1143 = _T_639 ? _T_284 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1145 = _T_641 ? _T_287 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1147 = _T_643 ? _T_287 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1149 = _T_645 ? _T_290 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1151 = _T_647 ? _T_290 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1153 = _T_649 ? _T_293 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1155 = _T_651 ? _T_293 : 40'h0; // @[Mux.scala 19:72]
  wire [63:0] _T_1160 = _T_991 | _T_993; // @[Mux.scala 19:72]
  wire [63:0] _GEN_154 = {{48'd0}, _T_995}; // @[Mux.scala 19:72]
  wire [63:0] _T_1161 = _T_1160 | _GEN_154; // @[Mux.scala 19:72]
  wire [63:0] _GEN_155 = {{55'd0}, _T_1001}; // @[Mux.scala 19:72]
  wire [63:0] _T_1164 = _T_1161 | _GEN_155; // @[Mux.scala 19:72]
  wire [63:0] _GEN_156 = {{29'd0}, _T_1003}; // @[Mux.scala 19:72]
  wire [63:0] _T_1165 = _T_1164 | _GEN_156; // @[Mux.scala 19:72]
  wire [63:0] _GEN_157 = {{55'd0}, _T_1005}; // @[Mux.scala 19:72]
  wire [63:0] _T_1166 = _T_1165 | _GEN_157; // @[Mux.scala 19:72]
  wire [63:0] _GEN_158 = {{48'd0}, _T_1007}; // @[Mux.scala 19:72]
  wire [63:0] _T_1167 = _T_1166 | _GEN_158; // @[Mux.scala 19:72]
  wire [63:0] _GEN_159 = {{48'd0}, _T_1009}; // @[Mux.scala 19:72]
  wire [63:0] _T_1168 = _T_1167 | _GEN_159; // @[Mux.scala 19:72]
  wire [63:0] _GEN_160 = {{32'd0}, _T_1011}; // @[Mux.scala 19:72]
  wire [63:0] _T_1169 = _T_1168 | _GEN_160; // @[Mux.scala 19:72]
  wire [63:0] _GEN_161 = {{32'd0}, _T_1013}; // @[Mux.scala 19:72]
  wire [63:0] _T_1170 = _T_1169 | _GEN_161; // @[Mux.scala 19:72]
  wire [63:0] _GEN_162 = {{32'd0}, _T_1015}; // @[Mux.scala 19:72]
  wire [63:0] _T_1171 = _T_1170 | _GEN_162; // @[Mux.scala 19:72]
  wire [63:0] _GEN_163 = {{32'd0}, _T_1017}; // @[Mux.scala 19:72]
  wire [63:0] _T_1172 = _T_1171 | _GEN_163; // @[Mux.scala 19:72]
  wire [63:0] _GEN_164 = {{32'd0}, _T_1021}; // @[Mux.scala 19:72]
  wire [63:0] _T_1174 = _T_1172 | _GEN_164; // @[Mux.scala 19:72]
  wire [63:0] _GEN_165 = {{32'd0}, _T_1023}; // @[Mux.scala 19:72]
  wire [63:0] _T_1175 = _T_1174 | _GEN_165; // @[Mux.scala 19:72]
  wire [63:0] _GEN_166 = {{32'd0}, _T_1025}; // @[Mux.scala 19:72]
  wire [63:0] _T_1176 = _T_1175 | _GEN_166; // @[Mux.scala 19:72]
  wire [63:0] _GEN_167 = {{32'd0}, _T_1027}; // @[Mux.scala 19:72]
  wire [63:0] _T_1177 = _T_1176 | _GEN_167; // @[Mux.scala 19:72]
  wire [63:0] _GEN_168 = {{24'd0}, _T_1029}; // @[Mux.scala 19:72]
  wire [63:0] _T_1178 = _T_1177 | _GEN_168; // @[Mux.scala 19:72]
  wire [63:0] _GEN_169 = {{24'd0}, _T_1031}; // @[Mux.scala 19:72]
  wire [63:0] _T_1179 = _T_1178 | _GEN_169; // @[Mux.scala 19:72]
  wire [63:0] _GEN_170 = {{24'd0}, _T_1033}; // @[Mux.scala 19:72]
  wire [63:0] _T_1180 = _T_1179 | _GEN_170; // @[Mux.scala 19:72]
  wire [63:0] _GEN_171 = {{24'd0}, _T_1035}; // @[Mux.scala 19:72]
  wire [63:0] _T_1181 = _T_1180 | _GEN_171; // @[Mux.scala 19:72]
  wire [63:0] _GEN_172 = {{24'd0}, _T_1037}; // @[Mux.scala 19:72]
  wire [63:0] _T_1182 = _T_1181 | _GEN_172; // @[Mux.scala 19:72]
  wire [63:0] _GEN_173 = {{24'd0}, _T_1039}; // @[Mux.scala 19:72]
  wire [63:0] _T_1183 = _T_1182 | _GEN_173; // @[Mux.scala 19:72]
  wire [63:0] _GEN_174 = {{24'd0}, _T_1041}; // @[Mux.scala 19:72]
  wire [63:0] _T_1184 = _T_1183 | _GEN_174; // @[Mux.scala 19:72]
  wire [63:0] _GEN_175 = {{24'd0}, _T_1043}; // @[Mux.scala 19:72]
  wire [63:0] _T_1185 = _T_1184 | _GEN_175; // @[Mux.scala 19:72]
  wire [63:0] _GEN_176 = {{24'd0}, _T_1045}; // @[Mux.scala 19:72]
  wire [63:0] _T_1186 = _T_1185 | _GEN_176; // @[Mux.scala 19:72]
  wire [63:0] _GEN_177 = {{24'd0}, _T_1047}; // @[Mux.scala 19:72]
  wire [63:0] _T_1187 = _T_1186 | _GEN_177; // @[Mux.scala 19:72]
  wire [63:0] _GEN_178 = {{24'd0}, _T_1049}; // @[Mux.scala 19:72]
  wire [63:0] _T_1188 = _T_1187 | _GEN_178; // @[Mux.scala 19:72]
  wire [63:0] _GEN_179 = {{24'd0}, _T_1051}; // @[Mux.scala 19:72]
  wire [63:0] _T_1189 = _T_1188 | _GEN_179; // @[Mux.scala 19:72]
  wire [63:0] _GEN_180 = {{24'd0}, _T_1053}; // @[Mux.scala 19:72]
  wire [63:0] _T_1190 = _T_1189 | _GEN_180; // @[Mux.scala 19:72]
  wire [63:0] _GEN_181 = {{24'd0}, _T_1055}; // @[Mux.scala 19:72]
  wire [63:0] _T_1191 = _T_1190 | _GEN_181; // @[Mux.scala 19:72]
  wire [63:0] _GEN_182 = {{24'd0}, _T_1057}; // @[Mux.scala 19:72]
  wire [63:0] _T_1192 = _T_1191 | _GEN_182; // @[Mux.scala 19:72]
  wire [63:0] _GEN_183 = {{24'd0}, _T_1059}; // @[Mux.scala 19:72]
  wire [63:0] _T_1193 = _T_1192 | _GEN_183; // @[Mux.scala 19:72]
  wire [63:0] _GEN_184 = {{24'd0}, _T_1061}; // @[Mux.scala 19:72]
  wire [63:0] _T_1194 = _T_1193 | _GEN_184; // @[Mux.scala 19:72]
  wire [63:0] _GEN_185 = {{24'd0}, _T_1063}; // @[Mux.scala 19:72]
  wire [63:0] _T_1195 = _T_1194 | _GEN_185; // @[Mux.scala 19:72]
  wire [63:0] _GEN_186 = {{24'd0}, _T_1065}; // @[Mux.scala 19:72]
  wire [63:0] _T_1196 = _T_1195 | _GEN_186; // @[Mux.scala 19:72]
  wire [63:0] _GEN_187 = {{24'd0}, _T_1067}; // @[Mux.scala 19:72]
  wire [63:0] _T_1197 = _T_1196 | _GEN_187; // @[Mux.scala 19:72]
  wire [63:0] _GEN_188 = {{24'd0}, _T_1069}; // @[Mux.scala 19:72]
  wire [63:0] _T_1198 = _T_1197 | _GEN_188; // @[Mux.scala 19:72]
  wire [63:0] _GEN_189 = {{24'd0}, _T_1071}; // @[Mux.scala 19:72]
  wire [63:0] _T_1199 = _T_1198 | _GEN_189; // @[Mux.scala 19:72]
  wire [63:0] _GEN_190 = {{24'd0}, _T_1073}; // @[Mux.scala 19:72]
  wire [63:0] _T_1200 = _T_1199 | _GEN_190; // @[Mux.scala 19:72]
  wire [63:0] _GEN_191 = {{24'd0}, _T_1075}; // @[Mux.scala 19:72]
  wire [63:0] _T_1201 = _T_1200 | _GEN_191; // @[Mux.scala 19:72]
  wire [63:0] _GEN_192 = {{24'd0}, _T_1077}; // @[Mux.scala 19:72]
  wire [63:0] _T_1202 = _T_1201 | _GEN_192; // @[Mux.scala 19:72]
  wire [63:0] _GEN_193 = {{24'd0}, _T_1079}; // @[Mux.scala 19:72]
  wire [63:0] _T_1203 = _T_1202 | _GEN_193; // @[Mux.scala 19:72]
  wire [63:0] _GEN_194 = {{24'd0}, _T_1081}; // @[Mux.scala 19:72]
  wire [63:0] _T_1204 = _T_1203 | _GEN_194; // @[Mux.scala 19:72]
  wire [63:0] _GEN_195 = {{24'd0}, _T_1083}; // @[Mux.scala 19:72]
  wire [63:0] _T_1205 = _T_1204 | _GEN_195; // @[Mux.scala 19:72]
  wire [63:0] _GEN_196 = {{24'd0}, _T_1085}; // @[Mux.scala 19:72]
  wire [63:0] _T_1206 = _T_1205 | _GEN_196; // @[Mux.scala 19:72]
  wire [63:0] _GEN_197 = {{24'd0}, _T_1087}; // @[Mux.scala 19:72]
  wire [63:0] _T_1207 = _T_1206 | _GEN_197; // @[Mux.scala 19:72]
  wire [63:0] _GEN_198 = {{24'd0}, _T_1089}; // @[Mux.scala 19:72]
  wire [63:0] _T_1208 = _T_1207 | _GEN_198; // @[Mux.scala 19:72]
  wire [63:0] _GEN_199 = {{24'd0}, _T_1091}; // @[Mux.scala 19:72]
  wire [63:0] _T_1209 = _T_1208 | _GEN_199; // @[Mux.scala 19:72]
  wire [63:0] _GEN_200 = {{24'd0}, _T_1093}; // @[Mux.scala 19:72]
  wire [63:0] _T_1210 = _T_1209 | _GEN_200; // @[Mux.scala 19:72]
  wire [63:0] _GEN_201 = {{24'd0}, _T_1095}; // @[Mux.scala 19:72]
  wire [63:0] _T_1211 = _T_1210 | _GEN_201; // @[Mux.scala 19:72]
  wire [63:0] _GEN_202 = {{24'd0}, _T_1097}; // @[Mux.scala 19:72]
  wire [63:0] _T_1212 = _T_1211 | _GEN_202; // @[Mux.scala 19:72]
  wire [63:0] _GEN_203 = {{24'd0}, _T_1099}; // @[Mux.scala 19:72]
  wire [63:0] _T_1213 = _T_1212 | _GEN_203; // @[Mux.scala 19:72]
  wire [63:0] _GEN_204 = {{24'd0}, _T_1101}; // @[Mux.scala 19:72]
  wire [63:0] _T_1214 = _T_1213 | _GEN_204; // @[Mux.scala 19:72]
  wire [63:0] _GEN_205 = {{24'd0}, _T_1103}; // @[Mux.scala 19:72]
  wire [63:0] _T_1215 = _T_1214 | _GEN_205; // @[Mux.scala 19:72]
  wire [63:0] _GEN_206 = {{24'd0}, _T_1105}; // @[Mux.scala 19:72]
  wire [63:0] _T_1216 = _T_1215 | _GEN_206; // @[Mux.scala 19:72]
  wire [63:0] _GEN_207 = {{24'd0}, _T_1107}; // @[Mux.scala 19:72]
  wire [63:0] _T_1217 = _T_1216 | _GEN_207; // @[Mux.scala 19:72]
  wire [63:0] _GEN_208 = {{24'd0}, _T_1109}; // @[Mux.scala 19:72]
  wire [63:0] _T_1218 = _T_1217 | _GEN_208; // @[Mux.scala 19:72]
  wire [63:0] _GEN_209 = {{24'd0}, _T_1111}; // @[Mux.scala 19:72]
  wire [63:0] _T_1219 = _T_1218 | _GEN_209; // @[Mux.scala 19:72]
  wire [63:0] _GEN_210 = {{24'd0}, _T_1113}; // @[Mux.scala 19:72]
  wire [63:0] _T_1220 = _T_1219 | _GEN_210; // @[Mux.scala 19:72]
  wire [63:0] _GEN_211 = {{24'd0}, _T_1115}; // @[Mux.scala 19:72]
  wire [63:0] _T_1221 = _T_1220 | _GEN_211; // @[Mux.scala 19:72]
  wire [63:0] _GEN_212 = {{24'd0}, _T_1117}; // @[Mux.scala 19:72]
  wire [63:0] _T_1222 = _T_1221 | _GEN_212; // @[Mux.scala 19:72]
  wire [63:0] _GEN_213 = {{24'd0}, _T_1119}; // @[Mux.scala 19:72]
  wire [63:0] _T_1223 = _T_1222 | _GEN_213; // @[Mux.scala 19:72]
  wire [63:0] _GEN_214 = {{24'd0}, _T_1121}; // @[Mux.scala 19:72]
  wire [63:0] _T_1224 = _T_1223 | _GEN_214; // @[Mux.scala 19:72]
  wire [63:0] _GEN_215 = {{24'd0}, _T_1123}; // @[Mux.scala 19:72]
  wire [63:0] _T_1225 = _T_1224 | _GEN_215; // @[Mux.scala 19:72]
  wire [63:0] _GEN_216 = {{24'd0}, _T_1125}; // @[Mux.scala 19:72]
  wire [63:0] _T_1226 = _T_1225 | _GEN_216; // @[Mux.scala 19:72]
  wire [63:0] _GEN_217 = {{24'd0}, _T_1127}; // @[Mux.scala 19:72]
  wire [63:0] _T_1227 = _T_1226 | _GEN_217; // @[Mux.scala 19:72]
  wire [63:0] _GEN_218 = {{24'd0}, _T_1129}; // @[Mux.scala 19:72]
  wire [63:0] _T_1228 = _T_1227 | _GEN_218; // @[Mux.scala 19:72]
  wire [63:0] _GEN_219 = {{24'd0}, _T_1131}; // @[Mux.scala 19:72]
  wire [63:0] _T_1229 = _T_1228 | _GEN_219; // @[Mux.scala 19:72]
  wire [63:0] _GEN_220 = {{24'd0}, _T_1133}; // @[Mux.scala 19:72]
  wire [63:0] _T_1230 = _T_1229 | _GEN_220; // @[Mux.scala 19:72]
  wire [63:0] _GEN_221 = {{24'd0}, _T_1135}; // @[Mux.scala 19:72]
  wire [63:0] _T_1231 = _T_1230 | _GEN_221; // @[Mux.scala 19:72]
  wire [63:0] _GEN_222 = {{24'd0}, _T_1137}; // @[Mux.scala 19:72]
  wire [63:0] _T_1232 = _T_1231 | _GEN_222; // @[Mux.scala 19:72]
  wire [63:0] _GEN_223 = {{24'd0}, _T_1139}; // @[Mux.scala 19:72]
  wire [63:0] _T_1233 = _T_1232 | _GEN_223; // @[Mux.scala 19:72]
  wire [63:0] _GEN_224 = {{24'd0}, _T_1141}; // @[Mux.scala 19:72]
  wire [63:0] _T_1234 = _T_1233 | _GEN_224; // @[Mux.scala 19:72]
  wire [63:0] _GEN_225 = {{24'd0}, _T_1143}; // @[Mux.scala 19:72]
  wire [63:0] _T_1235 = _T_1234 | _GEN_225; // @[Mux.scala 19:72]
  wire [63:0] _GEN_226 = {{24'd0}, _T_1145}; // @[Mux.scala 19:72]
  wire [63:0] _T_1236 = _T_1235 | _GEN_226; // @[Mux.scala 19:72]
  wire [63:0] _GEN_227 = {{24'd0}, _T_1147}; // @[Mux.scala 19:72]
  wire [63:0] _T_1237 = _T_1236 | _GEN_227; // @[Mux.scala 19:72]
  wire [63:0] _GEN_228 = {{24'd0}, _T_1149}; // @[Mux.scala 19:72]
  wire [63:0] _T_1238 = _T_1237 | _GEN_228; // @[Mux.scala 19:72]
  wire [63:0] _GEN_229 = {{24'd0}, _T_1151}; // @[Mux.scala 19:72]
  wire [63:0] _T_1239 = _T_1238 | _GEN_229; // @[Mux.scala 19:72]
  wire [63:0] _GEN_230 = {{24'd0}, _T_1153}; // @[Mux.scala 19:72]
  wire [63:0] _T_1240 = _T_1239 | _GEN_230; // @[Mux.scala 19:72]
  wire [63:0] _GEN_231 = {{24'd0}, _T_1155}; // @[Mux.scala 19:72]
  wire [63:0] _T_1241 = _T_1240 | _GEN_231; // @[Mux.scala 19:72]
  wire [34:0] _T_1270 = {{3'd0}, wdata};
  wire [39:0] _T_1338 = {wdata[7:0],_T_200[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_24 = _T_527 ? {{1'd0}, _T_1338} : _T_201; // @[csr.scala 386:29]
  wire [39:0] _T_1340 = {_T_200[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_25 = _T_525 ? {{1'd0}, _T_1340} : _GEN_24; // @[csr.scala 387:29]
  wire [39:0] _T_1343 = {wdata[7:0],_T_203[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_26 = _T_531 ? {{1'd0}, _T_1343} : _T_204; // @[csr.scala 386:29]
  wire [39:0] _T_1345 = {_T_203[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_27 = _T_529 ? {{1'd0}, _T_1345} : _GEN_26; // @[csr.scala 387:29]
  wire [39:0] _T_1348 = {wdata[7:0],_T_206[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_28 = _T_535 ? {{1'd0}, _T_1348} : _T_207; // @[csr.scala 386:29]
  wire [39:0] _T_1350 = {_T_206[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_29 = _T_533 ? {{1'd0}, _T_1350} : _GEN_28; // @[csr.scala 387:29]
  wire [39:0] _T_1353 = {wdata[7:0],_T_209[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_30 = _T_539 ? {{1'd0}, _T_1353} : _T_210; // @[csr.scala 386:29]
  wire [39:0] _T_1355 = {_T_209[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_31 = _T_537 ? {{1'd0}, _T_1355} : _GEN_30; // @[csr.scala 387:29]
  wire [39:0] _T_1358 = {wdata[7:0],_T_212[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_32 = _T_543 ? {{1'd0}, _T_1358} : _T_213; // @[csr.scala 386:29]
  wire [39:0] _T_1360 = {_T_212[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_33 = _T_541 ? {{1'd0}, _T_1360} : _GEN_32; // @[csr.scala 387:29]
  wire [39:0] _T_1363 = {wdata[7:0],_T_215[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_34 = _T_547 ? {{1'd0}, _T_1363} : _T_216; // @[csr.scala 386:29]
  wire [39:0] _T_1365 = {_T_215[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_35 = _T_545 ? {{1'd0}, _T_1365} : _GEN_34; // @[csr.scala 387:29]
  wire [39:0] _T_1368 = {wdata[7:0],_T_218[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_36 = _T_551 ? {{1'd0}, _T_1368} : _T_219; // @[csr.scala 386:29]
  wire [39:0] _T_1370 = {_T_218[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_37 = _T_549 ? {{1'd0}, _T_1370} : _GEN_36; // @[csr.scala 387:29]
  wire [39:0] _T_1373 = {wdata[7:0],_T_221[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_38 = _T_555 ? {{1'd0}, _T_1373} : _T_222; // @[csr.scala 386:29]
  wire [39:0] _T_1375 = {_T_221[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_39 = _T_553 ? {{1'd0}, _T_1375} : _GEN_38; // @[csr.scala 387:29]
  wire [39:0] _T_1378 = {wdata[7:0],_T_224[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_40 = _T_559 ? {{1'd0}, _T_1378} : _T_225; // @[csr.scala 386:29]
  wire [39:0] _T_1380 = {_T_224[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_41 = _T_557 ? {{1'd0}, _T_1380} : _GEN_40; // @[csr.scala 387:29]
  wire [39:0] _T_1383 = {wdata[7:0],_T_227[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_42 = _T_563 ? {{1'd0}, _T_1383} : _T_228; // @[csr.scala 386:29]
  wire [39:0] _T_1385 = {_T_227[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_43 = _T_561 ? {{1'd0}, _T_1385} : _GEN_42; // @[csr.scala 387:29]
  wire [39:0] _T_1388 = {wdata[7:0],_T_230[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_44 = _T_567 ? {{1'd0}, _T_1388} : _T_231; // @[csr.scala 386:29]
  wire [39:0] _T_1390 = {_T_230[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_45 = _T_565 ? {{1'd0}, _T_1390} : _GEN_44; // @[csr.scala 387:29]
  wire [39:0] _T_1393 = {wdata[7:0],_T_233[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_46 = _T_571 ? {{1'd0}, _T_1393} : _T_234; // @[csr.scala 386:29]
  wire [39:0] _T_1395 = {_T_233[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_47 = _T_569 ? {{1'd0}, _T_1395} : _GEN_46; // @[csr.scala 387:29]
  wire [39:0] _T_1398 = {wdata[7:0],_T_236[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_48 = _T_575 ? {{1'd0}, _T_1398} : _T_237; // @[csr.scala 386:29]
  wire [39:0] _T_1400 = {_T_236[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_49 = _T_573 ? {{1'd0}, _T_1400} : _GEN_48; // @[csr.scala 387:29]
  wire [39:0] _T_1403 = {wdata[7:0],_T_239[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_50 = _T_579 ? {{1'd0}, _T_1403} : _T_240; // @[csr.scala 386:29]
  wire [39:0] _T_1405 = {_T_239[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_51 = _T_577 ? {{1'd0}, _T_1405} : _GEN_50; // @[csr.scala 387:29]
  wire [39:0] _T_1408 = {wdata[7:0],_T_242[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_52 = _T_583 ? {{1'd0}, _T_1408} : _T_243; // @[csr.scala 386:29]
  wire [39:0] _T_1410 = {_T_242[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_53 = _T_581 ? {{1'd0}, _T_1410} : _GEN_52; // @[csr.scala 387:29]
  wire [39:0] _T_1413 = {wdata[7:0],_T_245[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_54 = _T_587 ? {{1'd0}, _T_1413} : _T_246; // @[csr.scala 386:29]
  wire [39:0] _T_1415 = {_T_245[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_55 = _T_585 ? {{1'd0}, _T_1415} : _GEN_54; // @[csr.scala 387:29]
  wire [39:0] _T_1418 = {wdata[7:0],_T_248[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_56 = _T_591 ? {{1'd0}, _T_1418} : _T_249; // @[csr.scala 386:29]
  wire [39:0] _T_1420 = {_T_248[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_57 = _T_589 ? {{1'd0}, _T_1420} : _GEN_56; // @[csr.scala 387:29]
  wire [39:0] _T_1423 = {wdata[7:0],_T_251[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_58 = _T_595 ? {{1'd0}, _T_1423} : _T_252; // @[csr.scala 386:29]
  wire [39:0] _T_1425 = {_T_251[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_59 = _T_593 ? {{1'd0}, _T_1425} : _GEN_58; // @[csr.scala 387:29]
  wire [39:0] _T_1428 = {wdata[7:0],_T_254[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_60 = _T_599 ? {{1'd0}, _T_1428} : _T_255; // @[csr.scala 386:29]
  wire [39:0] _T_1430 = {_T_254[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_61 = _T_597 ? {{1'd0}, _T_1430} : _GEN_60; // @[csr.scala 387:29]
  wire [39:0] _T_1433 = {wdata[7:0],_T_257[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_62 = _T_603 ? {{1'd0}, _T_1433} : _T_258; // @[csr.scala 386:29]
  wire [39:0] _T_1435 = {_T_257[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_63 = _T_601 ? {{1'd0}, _T_1435} : _GEN_62; // @[csr.scala 387:29]
  wire [39:0] _T_1438 = {wdata[7:0],_T_260[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_64 = _T_607 ? {{1'd0}, _T_1438} : _T_261; // @[csr.scala 386:29]
  wire [39:0] _T_1440 = {_T_260[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_65 = _T_605 ? {{1'd0}, _T_1440} : _GEN_64; // @[csr.scala 387:29]
  wire [39:0] _T_1443 = {wdata[7:0],_T_263[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_66 = _T_611 ? {{1'd0}, _T_1443} : _T_264; // @[csr.scala 386:29]
  wire [39:0] _T_1445 = {_T_263[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_67 = _T_609 ? {{1'd0}, _T_1445} : _GEN_66; // @[csr.scala 387:29]
  wire [39:0] _T_1448 = {wdata[7:0],_T_266[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_68 = _T_615 ? {{1'd0}, _T_1448} : _T_267; // @[csr.scala 386:29]
  wire [39:0] _T_1450 = {_T_266[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_69 = _T_613 ? {{1'd0}, _T_1450} : _GEN_68; // @[csr.scala 387:29]
  wire [39:0] _T_1453 = {wdata[7:0],_T_269[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_70 = _T_619 ? {{1'd0}, _T_1453} : _T_270; // @[csr.scala 386:29]
  wire [39:0] _T_1455 = {_T_269[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_71 = _T_617 ? {{1'd0}, _T_1455} : _GEN_70; // @[csr.scala 387:29]
  wire [39:0] _T_1458 = {wdata[7:0],_T_272[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_72 = _T_623 ? {{1'd0}, _T_1458} : _T_273; // @[csr.scala 386:29]
  wire [39:0] _T_1460 = {_T_272[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_73 = _T_621 ? {{1'd0}, _T_1460} : _GEN_72; // @[csr.scala 387:29]
  wire [39:0] _T_1463 = {wdata[7:0],_T_275[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_74 = _T_627 ? {{1'd0}, _T_1463} : _T_276; // @[csr.scala 386:29]
  wire [39:0] _T_1465 = {_T_275[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_75 = _T_625 ? {{1'd0}, _T_1465} : _GEN_74; // @[csr.scala 387:29]
  wire [39:0] _T_1468 = {wdata[7:0],_T_278[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_76 = _T_631 ? {{1'd0}, _T_1468} : _T_279; // @[csr.scala 386:29]
  wire [39:0] _T_1470 = {_T_278[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_77 = _T_629 ? {{1'd0}, _T_1470} : _GEN_76; // @[csr.scala 387:29]
  wire [39:0] _T_1473 = {wdata[7:0],_T_281[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_78 = _T_635 ? {{1'd0}, _T_1473} : _T_282; // @[csr.scala 386:29]
  wire [39:0] _T_1475 = {_T_281[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_79 = _T_633 ? {{1'd0}, _T_1475} : _GEN_78; // @[csr.scala 387:29]
  wire [39:0] _T_1478 = {wdata[7:0],_T_284[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_80 = _T_639 ? {{1'd0}, _T_1478} : _T_285; // @[csr.scala 386:29]
  wire [39:0] _T_1480 = {_T_284[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_81 = _T_637 ? {{1'd0}, _T_1480} : _GEN_80; // @[csr.scala 387:29]
  wire [39:0] _T_1483 = {wdata[7:0],_T_287[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_82 = _T_643 ? {{1'd0}, _T_1483} : _T_288; // @[csr.scala 386:29]
  wire [39:0] _T_1485 = {_T_287[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_83 = _T_641 ? {{1'd0}, _T_1485} : _GEN_82; // @[csr.scala 387:29]
  wire [39:0] _T_1488 = {wdata[7:0],_T_290[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_84 = _T_647 ? {{1'd0}, _T_1488} : _T_291; // @[csr.scala 386:29]
  wire [39:0] _T_1490 = {_T_290[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_85 = _T_645 ? {{1'd0}, _T_1490} : _GEN_84; // @[csr.scala 387:29]
  wire [39:0] _T_1493 = {wdata[7:0],_T_293[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_86 = _T_651 ? {{1'd0}, _T_1493} : _T_294; // @[csr.scala 386:29]
  wire [39:0] _T_1495 = {_T_293[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_87 = _T_649 ? {{1'd0}, _T_1495} : _GEN_86; // @[csr.scala 387:29]
  wire [63:0] _T_1498 = {wdata,_T_185[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_88 = _T_653 ? _T_1498 : {{57'd0}, _T_177}; // @[csr.scala 386:29]
  wire [63:0] _T_1501 = {_T_185[63:32],wdata}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_90 = _T_487 ? _T_1501 : _GEN_88; // @[csr.scala 387:29]
  wire [63:0] _T_1505 = {wdata,_T_197[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_92 = _T_655 ? _T_1505 : {{57'd0}, _T_189}; // @[csr.scala 386:29]
  wire [63:0] _T_1508 = {_T_197[63:32],wdata}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_94 = _T_489 ? _T_1508 : _GEN_92; // @[csr.scala 387:29]
  wire [31:0] _T_1512 = {{2'd0}, wdata[31:2]}; // @[csr.scala 368:78]
  wire [33:0] _GEN_233 = {_T_1512, 2'h0}; // @[csr.scala 368:86]
  wire [34:0] _T_1514 = {{1'd0}, _GEN_233}; // @[csr.scala 368:86]
  wire [34:0] _GEN_98 = _T_509 ? _T_1514 : {{3'd0}, _GEN_4}; // @[csr.scala 368:40]
  wire [31:0] _T_1516 = wdata & 32'h8000001f; // @[csr.scala 370:62]
  wire [40:0] _GEN_110 = wen ? _GEN_25 : _T_201; // @[csr.scala 331:14]
  wire [40:0] _GEN_111 = wen ? _GEN_27 : _T_204; // @[csr.scala 331:14]
  wire [40:0] _GEN_112 = wen ? _GEN_29 : _T_207; // @[csr.scala 331:14]
  wire [40:0] _GEN_113 = wen ? _GEN_31 : _T_210; // @[csr.scala 331:14]
  wire [40:0] _GEN_114 = wen ? _GEN_33 : _T_213; // @[csr.scala 331:14]
  wire [40:0] _GEN_115 = wen ? _GEN_35 : _T_216; // @[csr.scala 331:14]
  wire [40:0] _GEN_116 = wen ? _GEN_37 : _T_219; // @[csr.scala 331:14]
  wire [40:0] _GEN_117 = wen ? _GEN_39 : _T_222; // @[csr.scala 331:14]
  wire [40:0] _GEN_118 = wen ? _GEN_41 : _T_225; // @[csr.scala 331:14]
  wire [40:0] _GEN_119 = wen ? _GEN_43 : _T_228; // @[csr.scala 331:14]
  wire [40:0] _GEN_120 = wen ? _GEN_45 : _T_231; // @[csr.scala 331:14]
  wire [40:0] _GEN_121 = wen ? _GEN_47 : _T_234; // @[csr.scala 331:14]
  wire [40:0] _GEN_122 = wen ? _GEN_49 : _T_237; // @[csr.scala 331:14]
  wire [40:0] _GEN_123 = wen ? _GEN_51 : _T_240; // @[csr.scala 331:14]
  wire [40:0] _GEN_124 = wen ? _GEN_53 : _T_243; // @[csr.scala 331:14]
  wire [40:0] _GEN_125 = wen ? _GEN_55 : _T_246; // @[csr.scala 331:14]
  wire [40:0] _GEN_126 = wen ? _GEN_57 : _T_249; // @[csr.scala 331:14]
  wire [40:0] _GEN_127 = wen ? _GEN_59 : _T_252; // @[csr.scala 331:14]
  wire [40:0] _GEN_128 = wen ? _GEN_61 : _T_255; // @[csr.scala 331:14]
  wire [40:0] _GEN_129 = wen ? _GEN_63 : _T_258; // @[csr.scala 331:14]
  wire [40:0] _GEN_130 = wen ? _GEN_65 : _T_261; // @[csr.scala 331:14]
  wire [40:0] _GEN_131 = wen ? _GEN_67 : _T_264; // @[csr.scala 331:14]
  wire [40:0] _GEN_132 = wen ? _GEN_69 : _T_267; // @[csr.scala 331:14]
  wire [40:0] _GEN_133 = wen ? _GEN_71 : _T_270; // @[csr.scala 331:14]
  wire [40:0] _GEN_134 = wen ? _GEN_73 : _T_273; // @[csr.scala 331:14]
  wire [40:0] _GEN_135 = wen ? _GEN_75 : _T_276; // @[csr.scala 331:14]
  wire [40:0] _GEN_136 = wen ? _GEN_77 : _T_279; // @[csr.scala 331:14]
  wire [40:0] _GEN_137 = wen ? _GEN_79 : _T_282; // @[csr.scala 331:14]
  wire [40:0] _GEN_138 = wen ? _GEN_81 : _T_285; // @[csr.scala 331:14]
  wire [40:0] _GEN_139 = wen ? _GEN_83 : _T_288; // @[csr.scala 331:14]
  wire [40:0] _GEN_140 = wen ? _GEN_85 : _T_291; // @[csr.scala 331:14]
  wire [40:0] _GEN_141 = wen ? _GEN_87 : _T_294; // @[csr.scala 331:14]
  wire [63:0] _GEN_142 = wen ? _GEN_90 : {{57'd0}, _T_177}; // @[csr.scala 331:14]
  wire [63:0] _GEN_144 = wen ? _GEN_94 : {{57'd0}, _T_189}; // @[csr.scala 331:14]
  wire [34:0] _GEN_148 = wen ? _GEN_98 : {{3'd0}, _GEN_4}; // @[csr.scala 331:14]
  assign io_rw_rdata = _T_1241[31:0]; // @[csr.scala 329:15]
  assign io_eret = _T_962 | insn_ret; // @[csr.scala 282:11]
  assign io_status_debug = 1'h0; // @[csr.scala 280:13]
  assign io_status_prv = 2'h3; // @[csr.scala 280:13]
  assign io_status_sd = 1'h0; // @[csr.scala 280:13]
  assign io_status_zero1 = 8'h0; // @[csr.scala 280:13]
  assign io_status_tsr = 1'h0; // @[csr.scala 280:13]
  assign io_status_tw = 1'h0; // @[csr.scala 280:13]
  assign io_status_tvm = 1'h0; // @[csr.scala 280:13]
  assign io_status_mxr = 1'h0; // @[csr.scala 280:13]
  assign io_status_sum = 1'h0; // @[csr.scala 280:13]
  assign io_status_mprv = 1'h0; // @[csr.scala 280:13]
  assign io_status_xs = 2'h0; // @[csr.scala 280:13]
  assign io_status_fs = 2'h0; // @[csr.scala 280:13]
  assign io_status_mpp = 2'h3; // @[csr.scala 280:13]
  assign io_status_hpp = 2'h0; // @[csr.scala 280:13]
  assign io_status_spp = 1'h0; // @[csr.scala 280:13]
  assign io_status_mpie = reg_mstatus_mpie; // @[csr.scala 280:13]
  assign io_status_hpie = 1'h0; // @[csr.scala 280:13]
  assign io_status_spie = 1'h0; // @[csr.scala 280:13]
  assign io_status_upie = 1'h0; // @[csr.scala 280:13]
  assign io_status_mie = reg_mstatus_mie; // @[csr.scala 280:13]
  assign io_status_hie = 1'h0; // @[csr.scala 280:13]
  assign io_status_sie = 1'h0; // @[csr.scala 280:13]
  assign io_status_uie = 1'h0; // @[csr.scala 280:13]
  assign io_evec = insn_break ? 32'h80000004 : _GEN_13; // @[csr.scala 287:13 csr.scala 301:13 csr.scala 309:13 csr.scala 314:13 csr.scala 320:13]
  assign _GEN_451_0 = reset;
  assign _GEN_331_0 = io_decode_csr == 12'hb88;
  assign _GEN_337_0 = io_decode_csr == 12'hb8b;
  assign _GEN_415_0 = cpu_wen & _T_663;
  assign _GEN_436_0 = cpu_wen & _T_663;
  assign _GEN_352_0 = io_decode_csr == 12'hb12;
  assign _GEN_430_0 = cpu_wen & _T_663;
  assign _GEN_151_0 = system_insn & opcode[0];
  assign _GEN_310_0 = io_decode_csr == 12'hb21;
  assign _GEN_409_0 = cpu_wen & _T_663;
  assign _GEN_253_0 = io_decode_csr == 12'hb84;
  assign _GEN_316_0 = io_decode_csr == 12'h300;
  assign _GEN_244_0 = io_decode_csr == 12'h343;
  assign _GEN_238_0 = io_decode_csr == 12'h300;
  assign _GEN_325_0 = io_decode_csr == 12'hb85;
  assign _GEN_433_0 = cpu_wen & _T_663;
  assign _GEN_313_0 = io_decode_csr == 12'hba2;
  assign _GEN_11_0 = io_exception;
  assign _GEN_304_0 = io_decode_csr == 12'hb1e;
  assign _GEN_294_0 = io_decode_csr == 12'hb19;
  assign _GEN_303_0 = io_decode_csr == 12'hb9d;
  assign _GEN_402_0 = cpu_wen & _T_663;
  assign _GEN_412_0 = cpu_wen & _T_663;
  assign _GEN_424_0 = cpu_wen & _T_663;
  assign _GEN_319_0 = io_decode_csr == 12'h304;
  assign _GEN_288_0 = io_decode_csr == 12'hb16;
  assign _GEN_418_0 = cpu_wen & _T_663;
  assign _GEN_387_0 = io_decode_csr == 12'hb00;
  assign _GEN_462_0 = reset;
  assign _GEN_375_0 = io_decode_csr == 12'hb9e;
  assign _GEN_390_0 = io_decode_csr == 12'hb82;
  assign _GEN_307_0 = io_decode_csr == 12'hb9f;
  assign _GEN_297_0 = io_decode_csr == 12'hb9a;
  assign _GEN_406_0 = cpu_wen & _T_663;
  assign _GEN_270_0 = io_decode_csr == 12'hb0d;
  assign _GEN_369_0 = io_decode_csr == 12'hb9b;
  assign _GEN_396_0 = io_decode_csr == 12'h340;
  assign _GEN_276_0 = io_decode_csr == 12'hb10;
  assign _GEN_291_0 = io_decode_csr == 12'hb97;
  assign _GEN_258_0 = io_decode_csr == 12'hb07;
  assign _GEN_372_0 = io_decode_csr == 12'hb1c;
  assign _GEN_252_1 = io_decode_csr == 12'hb04;
  assign _GEN_285_0 = io_decode_csr == 12'hb94;
  assign _GEN_384_0 = io_decode_csr == 12'hb22;
  assign _GEN_378_0 = io_decode_csr == 12'hb1f;
  assign _GEN_393_0 = io_decode_csr == 12'h7b1;
  assign _GEN_273_0 = io_decode_csr == 12'hb8e;
  assign _GEN_456_0 = reset;
  assign _GEN_351_1 = io_decode_csr == 12'hb92;
  assign _GEN_450_0 = cpu_wen & _T_663;
  assign _GEN_357_0 = io_decode_csr == 12'hb95;
  assign _GEN_279_0 = io_decode_csr == 12'hb91;
  assign _GEN_399_0 = io_decode_csr == 12'h302;
  assign _GEN_264_0 = io_decode_csr == 12'hb0a;
  assign _GEN_300_0 = io_decode_csr == 12'hb1c;
  assign _GEN_432_0 = cpu_wen & _T_663;
  assign _GEN_381_0 = io_decode_csr == 12'hba1;
  assign _GEN_339_1 = io_decode_csr == 12'hb8c;
  assign _GEN_261_0 = io_decode_csr == 12'hb88;
  assign _GEN_360_0 = io_decode_csr == 12'hb16;
  assign _GEN_246_1 = io_decode_csr == 12'h7b0;
  assign _GEN_438_0 = cpu_wen & _T_663;
  assign _GEN_282_0 = io_decode_csr == 12'hb13;
  assign _GEN_345_1 = io_decode_csr == 12'hb8f;
  assign _GEN_240_1 = io_decode_csr == 12'h344;
  assign _GEN_444_0 = system_insn & opcode[1];
  assign _GEN_267_1 = io_decode_csr == 12'hb8b;
  assign _GEN_459_0 = cpu_wen & _T_663;
  assign _GEN_453_0 = reset;
  assign _GEN_366_0 = io_decode_csr == 12'hb19;
  assign _GEN_7_0 = io_rw_cmd == 3'h3;
  assign _GEN_324_1 = io_decode_csr == 12'hb04;
  assign _GEN_333_1 = io_decode_csr == 12'hb89;
  assign _GEN_342_0 = io_decode_csr == 12'hb0d;
  assign _GEN_405_0 = cpu_wen & _T_663;
  assign _GEN_420_1 = cpu_wen & _T_663;
  assign _GEN_306_0 = io_decode_csr == 12'hb1f;
  assign _GEN_3_0 = _T_177[6];
  assign _GEN_426_0 = cpu_wen & _T_663;
  assign _GEN_441_0 = cpu_wen & _T_663;
  assign _GEN_348_0 = io_decode_csr == 12'hb10;
  assign _GEN_255_0 = io_decode_csr == 12'hb85;
  assign _GEN_146_0 = insn_ret & io_decode_csr[10];
  assign _GEN_363_0 = io_decode_csr == 12'hb98;
  assign _GEN_321_1 = io_decode_csr == 12'hb83;
  assign _GEN_327_1 = io_decode_csr == 12'hb86;
  assign _GEN_354_0 = io_decode_csr == 12'hb13;
  assign _GEN_234_1 = io_decode_csr == 12'hb00;
  assign _GEN_249_1 = io_decode_csr == 12'h302;
  assign _GEN_243_0 = io_decode_csr == 12'h341;
  assign _GEN_447_0 = cpu_wen & _T_663;
  assign _GEN_330_1 = io_decode_csr == 12'hb07;
  assign _GEN_429_0 = cpu_wen & _T_663;
  assign _GEN_293_1 = io_decode_csr == 12'hb98;
  assign _GEN_414_1 = cpu_wen & _T_663;
  assign _GEN_309_0 = io_decode_csr == 12'hba0;
  assign _GEN_299_1 = io_decode_csr == 12'hb9b;
  assign _GEN_336_0 = io_decode_csr == 12'hb0a;
  assign _GEN_408_0 = cpu_wen & _T_663;
  assign _GEN_150_0 = system_insn & opcode[0];
  assign _GEN_435_0 = cpu_wen & _T_663;
  assign _GEN_392_1 = io_decode_csr == 12'hb02;
  assign _GEN_398_1 = io_decode_csr == 12'h343;
  assign _GEN_423_1 = cpu_wen & _T_663;
  assign _GEN_237_0 = io_decode_csr == 12'h301;
  assign _GEN_315_1 = io_decode_csr == 12'h7b0;
  assign _GEN_302_1 = io_decode_csr == 12'hb1d;
  assign _GEN_380_1 = io_decode_csr == 12'hb20;
  assign _GEN_318_1 = io_decode_csr == 12'h344;
  assign _GEN_287_1 = io_decode_csr == 12'hb95;
  assign _GEN_386_1 = io_decode_csr == 12'hb80;
  assign _GEN_281_1 = io_decode_csr == 12'hb92;
  assign _GEN_312_1 = io_decode_csr == 12'hb22;
  assign _GEN_417_1 = cpu_wen & _T_663;
  assign _GEN_411_1 = cpu_wen & _T_663;
  assign _GEN_401_1 = cpu_wen & _T_663;
  assign _GEN_374_1 = io_decode_csr == 12'hb1d;
  assign _GEN_368_1 = io_decode_csr == 12'hb1a;
  assign _GEN_383_1 = io_decode_csr == 12'hba2;
  assign _GEN_263_1 = io_decode_csr == 12'hb89;
  assign _GEN_446_0 = reset;
  assign _GEN_290_1 = io_decode_csr == 12'hb17;
  assign _GEN_389_1 = io_decode_csr == 12'hb82;
  assign _GEN_254_1 = io_decode_csr == 12'hb05;
  assign _GEN_461_0 = reset;
  assign _GEN_362_1 = io_decode_csr == 12'hb17;
  assign _GEN_296_1 = io_decode_csr == 12'hb1a;
  assign _GEN_395_1 = io_decode_csr == 12'h341;
  assign _GEN_275_1 = io_decode_csr == 12'hb8f;
  assign _GEN_269_1 = io_decode_csr == 12'hb8c;
  assign _GEN_278_1 = io_decode_csr == 12'hb11;
  assign _GEN_251_1 = io_decode_csr == 12'hb83;
  assign _GEN_455_0 = reset;
  assign _GEN_377_1 = io_decode_csr == 12'hb9f;
  assign _GEN_272_1 = io_decode_csr == 12'hb0e;
  assign _GEN_335_1 = io_decode_csr == 12'hb8a;
  assign _GEN_434_0 = cpu_wen & _T_663;
  assign _GEN_257_1 = io_decode_csr == 12'hb86;
  assign _GEN_443_0 = cpu_wen & _T_663;
  assign _GEN_356_1 = io_decode_csr == 12'hb14;
  assign _GEN_350_1 = io_decode_csr == 12'hb11;
  assign _GEN_428_0 = cpu_wen & _T_663;
  assign _GEN_449_0 = cpu_wen & _T_663;
  assign _GEN_236_1 = io_decode_csr == 12'hf13;
  assign _GEN_371_1 = io_decode_csr == 12'hb9c;
  assign _GEN_284_1 = io_decode_csr == 12'hb14;
  assign _GEN_416_1 = cpu_wen & _T_663;
  assign _GEN_260_1 = io_decode_csr == 12'hb08;
  assign _GEN_338_1 = io_decode_csr == 12'hb0b;
  assign _GEN_344_1 = io_decode_csr == 12'hb0e;
  assign _GEN_239_1 = io_decode_csr == 12'h305;
  assign _GEN_353_1 = io_decode_csr == 12'hb93;
  assign _GEN_266_1 = io_decode_csr == 12'hb0b;
  assign _GEN_452_0 = reset;
  assign _GEN_365_1 = io_decode_csr == 12'hb99;
  assign _GEN_6_0 = _T_664 | _T_665;
  assign _GEN_410_1 = cpu_wen & _T_663;
  assign _GEN_152_1 = system_insn & opcode[1];
  assign _GEN_437_0 = cpu_wen & _T_663;
  assign _GEN_332_1 = io_decode_csr == 12'hb08;
  assign _GEN_245_1 = io_decode_csr == 12'h342;
  assign _GEN_359_1 = io_decode_csr == 12'hb96;
  assign _GEN_431_0 = cpu_wen & _T_663;
  assign _GEN_458_0 = reset;
  assign _GEN_317_1 = io_decode_csr == 12'h300;
  assign _GEN_326_1 = io_decode_csr == 12'hb05;
  assign _GEN_341_1 = io_decode_csr == 12'hb8d;
  assign _GEN_394_1 = io_decode_csr == 12'h7b2;
  assign _GEN_248_1 = io_decode_csr == 12'h7b2;
  assign _GEN_347_1 = io_decode_csr == 12'hb90;
  assign _GEN_425_1 = cpu_wen & _T_663;
  assign _GEN_305_1 = io_decode_csr == 12'hb9e;
  assign _GEN_419_1 = cpu_wen & _T_663;
  assign _GEN_320_1 = io_decode_csr == 12'h304;
  assign _GEN_413_1 = cpu_wen & _T_663;
  assign _GEN_440_0 = cpu_wen & _T_663;
  assign _GEN_295_1 = io_decode_csr == 12'hb99;
  assign _GEN_404_1 = cpu_wen & _T_663;
  assign _GEN_403_1 = cpu_wen & _T_663;
  assign _GEN_242_1 = io_decode_csr == 12'h340;
  assign _GEN_15_1 = io_exception;
  assign _GEN_308_1 = io_decode_csr == 12'hb20;
  assign _GEN_149_1 = insn_ret & _T_980;
  assign _GEN_329_1 = io_decode_csr == 12'hb87;
  assign _GEN_292_1 = io_decode_csr == 12'hb18;
  assign _GEN_298_1 = io_decode_csr == 12'hb1b;
  assign _GEN_391_1 = io_decode_csr == 12'hb02;
  assign _GEN_314_1 = io_decode_csr == 12'h7b0;
  assign _GEN_323_1 = io_decode_csr == 12'hb84;
  assign _GEN_376_1 = io_decode_csr == 12'hb1e;
  assign _GEN_422_1 = cpu_wen & _T_663;
  assign _GEN_277_1 = io_decode_csr == 12'hb90;
  assign _GEN_407_1 = cpu_wen & _T_663;
  assign _GEN_397_1 = io_decode_csr == 12'h342;
  assign _GEN_379_1 = io_decode_csr == 12'hba0;
  assign _GEN_373_1 = io_decode_csr == 12'hb9d;
  assign _GEN_364_1 = io_decode_csr == 12'hb18;
  assign _GEN_259_1 = io_decode_csr == 12'hb87;
  assign _GEN_265_1 = io_decode_csr == 12'hb8a;
  assign _GEN_301_1 = io_decode_csr == 12'hb9c;
  assign _GEN_286_1 = io_decode_csr == 12'hb15;
  assign _GEN_400_1 = cpu_wen & _T_663;
  assign _GEN_358_1 = io_decode_csr == 12'hb15;
  assign _GEN_385_1 = io_decode_csr == 12'hb80;
  assign _GEN_457_0 = reset;
  assign _GEN_311_1 = io_decode_csr == 12'hba1;
  assign _GEN_280_1 = io_decode_csr == 12'hb12;
  assign _GEN_367_1 = io_decode_csr == 12'hb9a;
  assign _GEN_247_1 = io_decode_csr == 12'h7b1;
  assign _GEN_274_1 = io_decode_csr == 12'hb0f;
  assign _GEN_460_0 = cpu_wen & _T_663;
  assign _GEN_283_1 = io_decode_csr == 12'hb93;
  assign _GEN_388_1 = io_decode_csr == 12'hb00;
  assign _GEN_382_1 = io_decode_csr == 12'hb21;
  assign _GEN_268_1 = io_decode_csr == 12'hb0c;
  assign _GEN_346_1 = io_decode_csr == 12'hb0f;
  assign _GEN_340_1 = io_decode_csr == 12'hb0c;
  assign _GEN_439_0 = cpu_wen & _T_663;
  assign _GEN_262_1 = io_decode_csr == 12'hb09;
  assign _GEN_361_1 = io_decode_csr == 12'hb97;
  assign _GEN_241_1 = io_decode_csr == 12'h304;
  assign _GEN_445_0 = reset;
  assign _GEN_289_1 = io_decode_csr == 12'hb96;
  assign _GEN_421_1 = cpu_wen & _T_663;
  assign _GEN_427_0 = cpu_wen & _T_663;
  assign _GEN_454_0 = reset;
  assign _GEN_256_1 = io_decode_csr == 12'hb06;
  assign _GEN_5_2 = _T_189[6];
  assign _GEN_271_1 = io_decode_csr == 12'hb8d;
  assign _GEN_322_1 = io_decode_csr == 12'hb03;
  assign _GEN_334_1 = io_decode_csr == 12'hb09;
  assign _GEN_235_1 = io_decode_csr == 12'hb02;
  assign _GEN_349_1 = io_decode_csr == 12'hb91;
  assign _GEN_147_2 = insn_ret & _T_980;
  assign _GEN_448_0 = cpu_wen & _T_663;
  assign _GEN_442_0 = cpu_wen & _T_663;
  assign _GEN_343_1 = io_decode_csr == 12'hb8e;
  assign _GEN_355_1 = io_decode_csr == 12'hb94;
  assign _GEN_370_1 = io_decode_csr == 12'hb1b;
  assign _GEN_250_1 = io_decode_csr == 12'hb03;
  assign _GEN_463_0 = ~_T_970;
  assign _GEN_328_1 = io_decode_csr == 12'hb06;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mstatus_mpie = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_mstatus_mie = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  reg_mepc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_mcause = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_mtval = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_mscratch = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_medeleg = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_mip_mtip = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  reg_mip_msip = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  reg_mie_mtip = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  reg_mie_msip = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_176 = _RAND_11[5:0];
  _RAND_12 = {2{`RANDOM}};
  _T_180 = _RAND_12[57:0];
  _RAND_13 = {1{`RANDOM}};
  _T_188 = _RAND_13[5:0];
  _RAND_14 = {2{`RANDOM}};
  _T_192 = _RAND_14[57:0];
  _RAND_15 = {2{`RANDOM}};
  _T_200 = _RAND_15[39:0];
  _RAND_16 = {2{`RANDOM}};
  _T_203 = _RAND_16[39:0];
  _RAND_17 = {2{`RANDOM}};
  _T_206 = _RAND_17[39:0];
  _RAND_18 = {2{`RANDOM}};
  _T_209 = _RAND_18[39:0];
  _RAND_19 = {2{`RANDOM}};
  _T_212 = _RAND_19[39:0];
  _RAND_20 = {2{`RANDOM}};
  _T_215 = _RAND_20[39:0];
  _RAND_21 = {2{`RANDOM}};
  _T_218 = _RAND_21[39:0];
  _RAND_22 = {2{`RANDOM}};
  _T_221 = _RAND_22[39:0];
  _RAND_23 = {2{`RANDOM}};
  _T_224 = _RAND_23[39:0];
  _RAND_24 = {2{`RANDOM}};
  _T_227 = _RAND_24[39:0];
  _RAND_25 = {2{`RANDOM}};
  _T_230 = _RAND_25[39:0];
  _RAND_26 = {2{`RANDOM}};
  _T_233 = _RAND_26[39:0];
  _RAND_27 = {2{`RANDOM}};
  _T_236 = _RAND_27[39:0];
  _RAND_28 = {2{`RANDOM}};
  _T_239 = _RAND_28[39:0];
  _RAND_29 = {2{`RANDOM}};
  _T_242 = _RAND_29[39:0];
  _RAND_30 = {2{`RANDOM}};
  _T_245 = _RAND_30[39:0];
  _RAND_31 = {2{`RANDOM}};
  _T_248 = _RAND_31[39:0];
  _RAND_32 = {2{`RANDOM}};
  _T_251 = _RAND_32[39:0];
  _RAND_33 = {2{`RANDOM}};
  _T_254 = _RAND_33[39:0];
  _RAND_34 = {2{`RANDOM}};
  _T_257 = _RAND_34[39:0];
  _RAND_35 = {2{`RANDOM}};
  _T_260 = _RAND_35[39:0];
  _RAND_36 = {2{`RANDOM}};
  _T_263 = _RAND_36[39:0];
  _RAND_37 = {2{`RANDOM}};
  _T_266 = _RAND_37[39:0];
  _RAND_38 = {2{`RANDOM}};
  _T_269 = _RAND_38[39:0];
  _RAND_39 = {2{`RANDOM}};
  _T_272 = _RAND_39[39:0];
  _RAND_40 = {2{`RANDOM}};
  _T_275 = _RAND_40[39:0];
  _RAND_41 = {2{`RANDOM}};
  _T_278 = _RAND_41[39:0];
  _RAND_42 = {2{`RANDOM}};
  _T_281 = _RAND_42[39:0];
  _RAND_43 = {2{`RANDOM}};
  _T_284 = _RAND_43[39:0];
  _RAND_44 = {2{`RANDOM}};
  _T_287 = _RAND_44[39:0];
  _RAND_45 = {2{`RANDOM}};
  _T_290 = _RAND_45[39:0];
  _RAND_46 = {2{`RANDOM}};
  _T_293 = _RAND_46[39:0];
  _RAND_47 = {1{`RANDOM}};
  reg_dpc = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  reg_dscratch = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  reg_dcsr_ebreakm = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  reg_dcsr_step = _RAND_50[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      reg_mstatus_mpie <= 1'h0;
    end else if (reset) begin
      reg_mstatus_mpie <= 1'h0;
    end else if (wen) begin
      if (_T_499) begin
        reg_mstatus_mpie <= _T_1270[7];
      end else begin
        reg_mstatus_mpie <= _GEN_10;
      end
    end else begin
      reg_mstatus_mpie <= _GEN_10;
    end
    if (metaReset) begin
      reg_mstatus_mie <= 1'h0;
    end else if (reset) begin
      reg_mstatus_mie <= 1'h0;
    end else if (wen) begin
      if (_T_499) begin
        reg_mstatus_mie <= _T_1270[3];
      end else if (_T_981) begin
        reg_mstatus_mie <= reg_mstatus_mpie;
      end
    end else if (_T_981) begin
      reg_mstatus_mie <= reg_mstatus_mpie;
    end
    if (metaReset) begin
      reg_mepc <= 32'h0;
    end else begin
      reg_mepc <= _GEN_148[31:0];
    end
    if (metaReset) begin
      reg_mcause <= 32'h0;
    end else if (wen) begin
      if (_T_513) begin
        reg_mcause <= _T_1516;
      end else if (insn_break) begin
        reg_mcause <= 32'h3;
      end else if (insn_call) begin
        reg_mcause <= 32'hb;
      end else if (io_exception) begin
        reg_mcause <= 32'h2;
      end
    end else if (insn_break) begin
      reg_mcause <= 32'h3;
    end else if (insn_call) begin
      reg_mcause <= 32'hb;
    end else if (io_exception) begin
      reg_mcause <= 32'h2;
    end
    if (metaReset) begin
      reg_mtval <= 32'h0;
    end else if (wen) begin
      if (_T_511) begin
        reg_mtval <= wdata;
      end
    end
    if (metaReset) begin
      reg_mscratch <= 32'h0;
    end else if (wen) begin
      if (_T_507) begin
        reg_mscratch <= wdata;
      end
    end
    if (metaReset) begin
      reg_medeleg <= 32'h0;
    end else if (wen) begin
      if (_T_523) begin
        reg_medeleg <= wdata;
      end
    end
    if (metaReset) begin
      reg_mip_mtip <= 1'h0;
    end else if (reset) begin
      reg_mip_mtip <= 1'h0;
    end else begin
      reg_mip_mtip <= 1'h1;
    end
    if (metaReset) begin
      reg_mip_msip <= 1'h0;
    end else if (reset) begin
      reg_mip_msip <= 1'h0;
    end else if (wen) begin
      if (_T_503) begin
        reg_mip_msip <= wdata[3];
      end
    end
    if (metaReset) begin
      reg_mie_mtip <= 1'h0;
    end else if (reset) begin
      reg_mie_mtip <= 1'h0;
    end else if (wen) begin
      if (_T_505) begin
        reg_mie_mtip <= wdata[7];
      end
    end
    if (metaReset) begin
      reg_mie_msip <= 1'h0;
    end else if (reset) begin
      reg_mie_msip <= 1'h0;
    end else if (wen) begin
      if (_T_505) begin
        reg_mie_msip <= wdata[3];
      end
    end
    if (metaReset) begin
      _T_176 <= 6'h0;
    end else if (reset) begin
      _T_176 <= 6'h0;
    end else begin
      _T_176 <= _GEN_142[5:0];
    end
    if (metaReset) begin
      _T_180 <= 58'h0;
    end else if (reset) begin
      _T_180 <= 58'h0;
    end else if (wen) begin
      if (_T_487) begin
        _T_180 <= _T_1501[63:6];
      end else if (_T_653) begin
        _T_180 <= _T_1498[63:6];
      end else if (_T_177[6]) begin
        _T_180 <= _T_184;
      end
    end else if (_T_177[6]) begin
      _T_180 <= _T_184;
    end
    if (metaReset) begin
      _T_188 <= 6'h0;
    end else if (reset) begin
      _T_188 <= 6'h0;
    end else begin
      _T_188 <= _GEN_144[5:0];
    end
    if (metaReset) begin
      _T_192 <= 58'h0;
    end else if (reset) begin
      _T_192 <= 58'h0;
    end else if (wen) begin
      if (_T_489) begin
        _T_192 <= _T_1508[63:6];
      end else if (_T_655) begin
        _T_192 <= _T_1505[63:6];
      end else if (_T_189[6]) begin
        _T_192 <= _T_196;
      end
    end else if (_T_189[6]) begin
      _T_192 <= _T_196;
    end
    if (metaReset) begin
      _T_200 <= 40'h0;
    end else begin
      _T_200 <= _GEN_110[39:0];
    end
    if (metaReset) begin
      _T_203 <= 40'h0;
    end else begin
      _T_203 <= _GEN_111[39:0];
    end
    if (metaReset) begin
      _T_206 <= 40'h0;
    end else begin
      _T_206 <= _GEN_112[39:0];
    end
    if (metaReset) begin
      _T_209 <= 40'h0;
    end else begin
      _T_209 <= _GEN_113[39:0];
    end
    if (metaReset) begin
      _T_212 <= 40'h0;
    end else begin
      _T_212 <= _GEN_114[39:0];
    end
    if (metaReset) begin
      _T_215 <= 40'h0;
    end else begin
      _T_215 <= _GEN_115[39:0];
    end
    if (metaReset) begin
      _T_218 <= 40'h0;
    end else begin
      _T_218 <= _GEN_116[39:0];
    end
    if (metaReset) begin
      _T_221 <= 40'h0;
    end else begin
      _T_221 <= _GEN_117[39:0];
    end
    if (metaReset) begin
      _T_224 <= 40'h0;
    end else begin
      _T_224 <= _GEN_118[39:0];
    end
    if (metaReset) begin
      _T_227 <= 40'h0;
    end else begin
      _T_227 <= _GEN_119[39:0];
    end
    if (metaReset) begin
      _T_230 <= 40'h0;
    end else begin
      _T_230 <= _GEN_120[39:0];
    end
    if (metaReset) begin
      _T_233 <= 40'h0;
    end else begin
      _T_233 <= _GEN_121[39:0];
    end
    if (metaReset) begin
      _T_236 <= 40'h0;
    end else begin
      _T_236 <= _GEN_122[39:0];
    end
    if (metaReset) begin
      _T_239 <= 40'h0;
    end else begin
      _T_239 <= _GEN_123[39:0];
    end
    if (metaReset) begin
      _T_242 <= 40'h0;
    end else begin
      _T_242 <= _GEN_124[39:0];
    end
    if (metaReset) begin
      _T_245 <= 40'h0;
    end else begin
      _T_245 <= _GEN_125[39:0];
    end
    if (metaReset) begin
      _T_248 <= 40'h0;
    end else begin
      _T_248 <= _GEN_126[39:0];
    end
    if (metaReset) begin
      _T_251 <= 40'h0;
    end else begin
      _T_251 <= _GEN_127[39:0];
    end
    if (metaReset) begin
      _T_254 <= 40'h0;
    end else begin
      _T_254 <= _GEN_128[39:0];
    end
    if (metaReset) begin
      _T_257 <= 40'h0;
    end else begin
      _T_257 <= _GEN_129[39:0];
    end
    if (metaReset) begin
      _T_260 <= 40'h0;
    end else begin
      _T_260 <= _GEN_130[39:0];
    end
    if (metaReset) begin
      _T_263 <= 40'h0;
    end else begin
      _T_263 <= _GEN_131[39:0];
    end
    if (metaReset) begin
      _T_266 <= 40'h0;
    end else begin
      _T_266 <= _GEN_132[39:0];
    end
    if (metaReset) begin
      _T_269 <= 40'h0;
    end else begin
      _T_269 <= _GEN_133[39:0];
    end
    if (metaReset) begin
      _T_272 <= 40'h0;
    end else begin
      _T_272 <= _GEN_134[39:0];
    end
    if (metaReset) begin
      _T_275 <= 40'h0;
    end else begin
      _T_275 <= _GEN_135[39:0];
    end
    if (metaReset) begin
      _T_278 <= 40'h0;
    end else begin
      _T_278 <= _GEN_136[39:0];
    end
    if (metaReset) begin
      _T_281 <= 40'h0;
    end else begin
      _T_281 <= _GEN_137[39:0];
    end
    if (metaReset) begin
      _T_284 <= 40'h0;
    end else begin
      _T_284 <= _GEN_138[39:0];
    end
    if (metaReset) begin
      _T_287 <= 40'h0;
    end else begin
      _T_287 <= _GEN_139[39:0];
    end
    if (metaReset) begin
      _T_290 <= 40'h0;
    end else begin
      _T_290 <= _GEN_140[39:0];
    end
    if (metaReset) begin
      _T_293 <= 40'h0;
    end else begin
      _T_293 <= _GEN_141[39:0];
    end
    if (metaReset) begin
      reg_dpc <= 32'h0;
    end else if (wen) begin
      if (_T_519) begin
        reg_dpc <= wdata;
      end
    end
    if (metaReset) begin
      reg_dscratch <= 32'h0;
    end else if (wen) begin
      if (_T_521) begin
        reg_dscratch <= wdata;
      end
    end
    if (metaReset) begin
      reg_dcsr_ebreakm <= 1'h0;
    end else if (reset) begin
      reg_dcsr_ebreakm <= 1'h0;
    end else if (wen) begin
      if (_T_517) begin
        reg_dcsr_ebreakm <= wdata[15];
      end
    end
    if (metaReset) begin
      reg_dcsr_step <= 1'h0;
    end else if (reset) begin
      reg_dcsr_step <= 1'h0;
    end else if (wen) begin
      if (_T_517) begin
        reg_dcsr_step <= wdata[2];
      end
    end
  end
endmodule
module DatPath(
  input         metaReset,
  input         clock,
  input         reset,
  output [31:0] io_imem_req_bits_addr,
  input  [31:0] io_imem_resp_bits_data,
  output        io_dmem_req_valid,
  output [31:0] io_dmem_req_bits_addr,
  output [31:0] io_dmem_req_bits_data,
  output        io_dmem_req_bits_fcn,
  output [2:0]  io_dmem_req_bits_typ,
  input  [31:0] io_dmem_resp_bits_data,
  input         io_ctl_dec_stall,
  input         io_ctl_full_stall,
  input  [1:0]  io_ctl_exe_pc_sel,
  input  [3:0]  io_ctl_br_type,
  input         io_ctl_if_kill,
  input         io_ctl_dec_kill,
  input  [1:0]  io_ctl_op1_sel,
  input  [2:0]  io_ctl_op2_sel,
  input  [3:0]  io_ctl_alu_fun,
  input  [1:0]  io_ctl_wb_sel,
  input         io_ctl_rf_wen,
  input         io_ctl_mem_val,
  input  [1:0]  io_ctl_mem_fcn,
  input  [2:0]  io_ctl_mem_typ,
  input  [2:0]  io_ctl_csr_cmd,
  input         io_ctl_fencei,
  input         io_ctl_pipeline_kill,
  input         io_ctl_mem_exception,
  output [31:0] io_dat_dec_inst,
  output        io_dat_exe_br_eq,
  output        io_dat_exe_br_lt,
  output        io_dat_exe_br_ltu,
  output [3:0]  io_dat_exe_br_type,
  output        io_dat_mem_ctrl_dmem_val,
  output        io_dat_csr_eret,
  output        _GEN_451,
  output        _GEN_331,
  output        _GEN_337,
  output        _GEN_113_0,
  output        _GEN_415,
  output        _GEN_436,
  output        _GEN_140_0,
  output        _GEN_98_0,
  output        _GEN_352,
  output        _GEN_125_0,
  output        _GEN_430,
  output        _GEN_119_0,
  output        _GEN_88_0,
  output        _GEN_151_0,
  output        _GEN_310,
  output        _GEN_104_0,
  output        _GEN_409,
  output        _GEN_253,
  output        _GEN_316,
  output        _GEN_244,
  output        _GEN_238,
  output        _GEN_101_0,
  output        _GEN_325,
  output        _GEN_169_0,
  output        _GEN_433,
  output        _GEN_313,
  output        _GEN_91_0,
  output        _GEN_11_0,
  output        _GEN_304,
  output        _GEN_294,
  output        _GEN_303,
  output        _GEN_107_0,
  output        _GEN_0_0,
  output        _GEN_402,
  output        _GEN_412,
  output        _GEN_424,
  output        _GEN_175_0,
  output        _GEN_319,
  output        _GEN_288,
  output        _GEN_56_0,
  output        _GEN_418,
  output        _GEN_122_0,
  output        _GEN_387,
  output        _GEN_72_0,
  output        _GEN_75_0,
  output        _GEN_85_0,
  output        _GEN_178_0,
  output        _GEN_157_0,
  output        _GEN_462,
  output        _GEN_69_0,
  output        _GEN_375,
  output        _GEN_151_1,
  output        _GEN_33_0,
  output        _GEN_390,
  output        _GEN_307,
  output        _GEN_297,
  output        _GEN_406,
  output        _GEN_270,
  output        _GEN_95_0,
  output        _GEN_45_0,
  output        _GEN_369,
  output        _GEN_396,
  output        _GEN_172_0,
  output        _GEN_276,
  output        _GEN_291,
  output        _GEN_258,
  output        _GEN_372,
  output        _GEN_252_0,
  output        _GEN_166_0,
  output        _GEN_285,
  output        _GEN_42_0,
  output        _GEN_384,
  output        _GEN_378,
  output        _GEN_393,
  output        _GEN_273,
  output        _GEN_456,
  output        _GEN_80_0,
  output        _GEN_351_0,
  output        _GEN_139_0,
  output        _GEN_145_0,
  output        _GEN_450,
  output        _GEN_53_1,
  output        _GEN_357,
  output        _GEN_160_0,
  output        _GEN_279,
  output        _GEN_133_0,
  output        _GEN_399,
  output        _GEN_264,
  output        _GEN_300,
  output        _GEN_127_0,
  output        _GEN_432,
  output        _GEN_381,
  output        _GEN_339_0,
  output        _GEN_261,
  output        _GEN_16_0,
  output        _GEN_360,
  output        _GEN_163_0,
  output        _GEN_246_0,
  output        _GEN_438,
  output        _GEN_282,
  output        _GEN_345_0,
  output        _GEN_121_0,
  output        _GEN_240_0,
  output        _GEN_148_0,
  output        _GEN_154_0,
  output        _GEN_444,
  output        _GEN_267_0,
  output        _GEN_459,
  output        _GEN_453,
  output        _GEN_366,
  output        _GEN_7_0,
  output        _GEN_142_0,
  output        _GEN_324_0,
  output        _GEN_333_0,
  output        _GEN_342,
  output        _GEN_405,
  output        _GEN_420_0,
  output        _GEN_306,
  output        _GEN_109_1,
  output        _GEN_103_0,
  output        _GEN_3_0,
  output        _GEN_136_0,
  output        _GEN_426,
  output        _GEN_441,
  output        _GEN_94_1,
  output        _GEN_348,
  output        _GEN_255,
  output        _GEN_115_0,
  output        _GEN_146_0,
  output        _GEN_363,
  output        _GEN_321_0,
  output        _GEN_327_0,
  output        _GEN_354,
  output        _GEN_234_0,
  output        _GEN_130_0,
  output        _GEN_249_0,
  output        _GEN_243,
  output        _GEN_447,
  output        _GEN_330_0,
  output        _GEN_429,
  output        _GEN_293_0,
  output        _GEN_87_0,
  output        _GEN_414_0,
  output        _GEN_309,
  output        _GEN_299_0,
  output        _GEN_336,
  output        _GEN_408,
  output        _GEN_112_0,
  output        _GEN_150_0,
  output        _GEN_435,
  output        _GEN_97_1,
  output        _GEN_124_0,
  output        _GEN_118_0,
  output        _GEN_392_0,
  output        _GEN_398_0,
  output        _GEN_423_0,
  output        _GEN_237,
  output        _GEN_315_0,
  output        _GEN_79_0,
  output        _GEN_1_2,
  output        _GEN_90_0,
  output        _GEN_162_0,
  output        _GEN_302_0,
  output        _GEN_106_1,
  output        _GEN_71_1,
  output        _GEN_380_0,
  output        _GEN_174_0,
  output        _GEN_318_0,
  output        _GEN_287_0,
  output        _GEN_386_0,
  output        _GEN_281_0,
  output        _GEN_312_0,
  output        _GEN_417_0,
  output        _GEN_411_0,
  output        _GEN_55_1,
  output        _GEN_100_1,
  output        _GEN_168_1,
  output        _GEN_401_0,
  output        _GEN_44_1,
  output        _GEN_74_1,
  output        _GEN_374_0,
  output        _GEN_368_0,
  output        _GEN_383_0,
  output        _GEN_263_0,
  output        _GEN_177_0,
  output        _GEN_171_0,
  output        _GEN_446,
  output        _GEN_290_0,
  output        _GEN_83_0,
  output        _GEN_135_1,
  output        _GEN_389_0,
  output        _GEN_93_0,
  output        _GEN_254_0,
  output        _GEN_21_0,
  output        _GEN_461,
  output        _GEN_362_0,
  output        _GEN_156_0,
  output        _GEN_150_1,
  output        _GEN_68_1,
  output        _GEN_296_0,
  output        _GEN_395_0,
  output        _GEN_275_0,
  output        _GEN_269_0,
  output        _GEN_278_0,
  output        _GEN_138_0,
  output        _GEN_251_0,
  output        _GEN_455,
  output        _GEN_377_0,
  output        _GEN_153_1,
  output        _GEN_272_0,
  output        _GEN_47_1,
  output        _GEN_335_0,
  output        _GEN_41_1,
  output        _GEN_434,
  output        _GEN_257_0,
  output        _GEN_443,
  output        _GEN_356_0,
  output        _GEN_350_0,
  output        _GEN_132_1,
  output        _GEN_144_0,
  output        _GEN_159_0,
  output        _GEN_428,
  output        _GEN_449,
  output        _GEN_117_1,
  output        _GEN_236_0,
  output        _GEN_371_0,
  output        _GEN_165_0,
  output        _GEN_284_0,
  output        _GEN_147_1,
  output        _GEN_416_0,
  output        _GEN_260_0,
  output        _GEN_105_1,
  output        _GEN_338_0,
  output        _GEN_141_1,
  output        _GEN_99_1,
  output        _GEN_344_0,
  output        _GEN_239_0,
  output        _GEN_353_0,
  output        _GEN_266_0,
  output        _GEN_452,
  output        _GEN_120_1,
  output        _GEN_365_0,
  output        _GEN_6_0,
  output        _GEN_410_0,
  output        _GEN_152_1,
  output        _GEN_437,
  output        _GEN_332_0,
  output        _GEN_126_1,
  output        _GEN_245_0,
  output        _GEN_359_0,
  output        _GEN_431,
  output        _GEN_458,
  output        _GEN_317_0,
  output        _GEN_326_0,
  output        _GEN_341_0,
  output        _GEN_1_3,
  output        _GEN_394_0,
  output        _GEN_248_0,
  output        _GEN_347_0,
  output        _GEN_92_1,
  output        _GEN_102_1,
  output        _GEN_425_0,
  output        _GEN_305_0,
  output        _GEN_419_0,
  output        _GEN_320_0,
  output        _GEN_108_1,
  output        _GEN_114_1,
  output        _GEN_123_1,
  output        _GEN_413_0,
  output        _GEN_440,
  output        _GEN_295_0,
  output        _GEN_129_1,
  output        _GEN_404_0,
  output        _GEN_403_0,
  output        _GEN_242_0,
  output        _GEN_15_1,
  output        _GEN_96_1,
  output        _GEN_86_1,
  output        _GEN_164_1,
  output        _GEN_308_0,
  output        _GEN_149_1,
  output        _GEN_329_0,
  output        _GEN_292_0,
  output        _GEN_298_0,
  output        _GEN_391_0,
  output        _GEN_314_0,
  output        _GEN_323_0,
  output        _GEN_376_0,
  output        _GEN_422_0,
  output        _GEN_277_0,
  output        _GEN_46_1,
  output        _GEN_111_1,
  output        _GEN_78_1,
  output        _GEN_407_0,
  output        _GEN_179_1,
  output        _GEN_397_0,
  output        _GEN_173_1,
  output        _GEN_70_1,
  output        _GEN_379_0,
  output        _GEN_82_1,
  output        _GEN_373_0,
  output        _GEN_54_1,
  output        _GEN_364_0,
  output        _GEN_259_0,
  output        _GEN_167_1,
  output        _GEN_43_1,
  output        _GEN_161_1,
  output        _GEN_265_0,
  output        _GEN_301_0,
  output        _GEN_146_2,
  output        _GEN_286_0,
  output        _GEN_400_0,
  output        _GEN_89_0,
  output        _GEN_358_0,
  output        _GEN_385_0,
  output        _GEN_457,
  output        _GEN_311_0,
  output        _GEN_280_0,
  output        _GEN_143_1,
  output        _GEN_367_0,
  output        _GEN_247_0,
  output        _GEN_274_0,
  output        _GEN_460,
  output        _GEN_283_0,
  output        _GEN_388_0,
  output        _GEN_382_0,
  output        _GEN_268_0,
  output        _GEN_176_1,
  output        _GEN_346_0,
  output        _GEN_64_1,
  output        _GEN_340_0,
  output        _GEN_134_1,
  output        _GEN_149_2,
  output        _GEN_439,
  output        _GEN_262_0,
  output        _GEN_17_1,
  output        _GEN_361_0,
  output        _GEN_155_1,
  output        _GEN_170_1,
  output        _GEN_73_1,
  output        _GEN_128_1,
  output        _GEN_241_0,
  output        _GEN_445,
  output        _GEN_289_0,
  output        _GEN_131_1,
  output        _GEN_152_2,
  output        _GEN_421_0,
  output        _GEN_427,
  output        _GEN_454,
  output        _GEN_256_0,
  output        _GEN_110_1,
  output        _GEN_40_1,
  output        _GEN_5_2,
  output        _GEN_158_1,
  output        _GEN_271_0,
  output        _GEN_322_0,
  output        _GEN_334_0,
  output        _GEN_116_1,
  output        _GEN_235_0,
  output        _GEN_349_0,
  output        _GEN_147_2,
  output        _GEN_448,
  output        _GEN_442,
  output        _GEN_343_0,
  output        _GEN_355_0,
  output        _GEN_137_1,
  output        _GEN_370_0,
  output        _GEN_250_0,
  output        _GEN_463,
  output        _GEN_328_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire  regfile_metaReset; // @[dpath.scala 157:24]
  wire  regfile_clock; // @[dpath.scala 157:24]
  wire [4:0] regfile_io_rs1_addr; // @[dpath.scala 157:24]
  wire [31:0] regfile_io_rs1_data; // @[dpath.scala 157:24]
  wire [4:0] regfile_io_rs2_addr; // @[dpath.scala 157:24]
  wire [31:0] regfile_io_rs2_data; // @[dpath.scala 157:24]
  wire [4:0] regfile_io_waddr; // @[dpath.scala 157:24]
  wire [31:0] regfile_io_wdata; // @[dpath.scala 157:24]
  wire  regfile_io_wen; // @[dpath.scala 157:24]
  wire  regfile__GEN_0_0; // @[dpath.scala 157:24]
  wire  regfile__GEN_1_3; // @[dpath.scala 157:24]
  wire  csr_metaReset; // @[dpath.scala 356:20]
  wire  csr_clock; // @[dpath.scala 356:20]
  wire  csr_reset; // @[dpath.scala 356:20]
  wire [2:0] csr_io_rw_cmd; // @[dpath.scala 356:20]
  wire [31:0] csr_io_rw_rdata; // @[dpath.scala 356:20]
  wire [31:0] csr_io_rw_wdata; // @[dpath.scala 356:20]
  wire  csr_io_eret; // @[dpath.scala 356:20]
  wire [11:0] csr_io_decode_csr; // @[dpath.scala 356:20]
  wire  csr_io_status_debug; // @[dpath.scala 356:20]
  wire [1:0] csr_io_status_prv; // @[dpath.scala 356:20]
  wire  csr_io_status_sd; // @[dpath.scala 356:20]
  wire [7:0] csr_io_status_zero1; // @[dpath.scala 356:20]
  wire  csr_io_status_tsr; // @[dpath.scala 356:20]
  wire  csr_io_status_tw; // @[dpath.scala 356:20]
  wire  csr_io_status_tvm; // @[dpath.scala 356:20]
  wire  csr_io_status_mxr; // @[dpath.scala 356:20]
  wire  csr_io_status_sum; // @[dpath.scala 356:20]
  wire  csr_io_status_mprv; // @[dpath.scala 356:20]
  wire [1:0] csr_io_status_xs; // @[dpath.scala 356:20]
  wire [1:0] csr_io_status_fs; // @[dpath.scala 356:20]
  wire [1:0] csr_io_status_mpp; // @[dpath.scala 356:20]
  wire [1:0] csr_io_status_hpp; // @[dpath.scala 356:20]
  wire  csr_io_status_spp; // @[dpath.scala 356:20]
  wire  csr_io_status_mpie; // @[dpath.scala 356:20]
  wire  csr_io_status_hpie; // @[dpath.scala 356:20]
  wire  csr_io_status_spie; // @[dpath.scala 356:20]
  wire  csr_io_status_upie; // @[dpath.scala 356:20]
  wire  csr_io_status_mie; // @[dpath.scala 356:20]
  wire  csr_io_status_hie; // @[dpath.scala 356:20]
  wire  csr_io_status_sie; // @[dpath.scala 356:20]
  wire  csr_io_status_uie; // @[dpath.scala 356:20]
  wire [31:0] csr_io_evec; // @[dpath.scala 356:20]
  wire  csr_io_exception; // @[dpath.scala 356:20]
  wire  csr_io_retire; // @[dpath.scala 356:20]
  wire [31:0] csr_io_pc; // @[dpath.scala 356:20]
  wire  csr__GEN_451_0; // @[dpath.scala 356:20]
  wire  csr__GEN_331_0; // @[dpath.scala 356:20]
  wire  csr__GEN_337_0; // @[dpath.scala 356:20]
  wire  csr__GEN_415_0; // @[dpath.scala 356:20]
  wire  csr__GEN_436_0; // @[dpath.scala 356:20]
  wire  csr__GEN_352_0; // @[dpath.scala 356:20]
  wire  csr__GEN_430_0; // @[dpath.scala 356:20]
  wire  csr__GEN_151_0; // @[dpath.scala 356:20]
  wire  csr__GEN_310_0; // @[dpath.scala 356:20]
  wire  csr__GEN_409_0; // @[dpath.scala 356:20]
  wire  csr__GEN_253_0; // @[dpath.scala 356:20]
  wire  csr__GEN_316_0; // @[dpath.scala 356:20]
  wire  csr__GEN_244_0; // @[dpath.scala 356:20]
  wire  csr__GEN_238_0; // @[dpath.scala 356:20]
  wire  csr__GEN_325_0; // @[dpath.scala 356:20]
  wire  csr__GEN_433_0; // @[dpath.scala 356:20]
  wire  csr__GEN_313_0; // @[dpath.scala 356:20]
  wire  csr__GEN_11_0; // @[dpath.scala 356:20]
  wire  csr__GEN_304_0; // @[dpath.scala 356:20]
  wire  csr__GEN_294_0; // @[dpath.scala 356:20]
  wire  csr__GEN_303_0; // @[dpath.scala 356:20]
  wire  csr__GEN_402_0; // @[dpath.scala 356:20]
  wire  csr__GEN_412_0; // @[dpath.scala 356:20]
  wire  csr__GEN_424_0; // @[dpath.scala 356:20]
  wire  csr__GEN_319_0; // @[dpath.scala 356:20]
  wire  csr__GEN_288_0; // @[dpath.scala 356:20]
  wire  csr__GEN_418_0; // @[dpath.scala 356:20]
  wire  csr__GEN_387_0; // @[dpath.scala 356:20]
  wire  csr__GEN_462_0; // @[dpath.scala 356:20]
  wire  csr__GEN_375_0; // @[dpath.scala 356:20]
  wire  csr__GEN_390_0; // @[dpath.scala 356:20]
  wire  csr__GEN_307_0; // @[dpath.scala 356:20]
  wire  csr__GEN_297_0; // @[dpath.scala 356:20]
  wire  csr__GEN_406_0; // @[dpath.scala 356:20]
  wire  csr__GEN_270_0; // @[dpath.scala 356:20]
  wire  csr__GEN_369_0; // @[dpath.scala 356:20]
  wire  csr__GEN_396_0; // @[dpath.scala 356:20]
  wire  csr__GEN_276_0; // @[dpath.scala 356:20]
  wire  csr__GEN_291_0; // @[dpath.scala 356:20]
  wire  csr__GEN_258_0; // @[dpath.scala 356:20]
  wire  csr__GEN_372_0; // @[dpath.scala 356:20]
  wire  csr__GEN_252_1; // @[dpath.scala 356:20]
  wire  csr__GEN_285_0; // @[dpath.scala 356:20]
  wire  csr__GEN_384_0; // @[dpath.scala 356:20]
  wire  csr__GEN_378_0; // @[dpath.scala 356:20]
  wire  csr__GEN_393_0; // @[dpath.scala 356:20]
  wire  csr__GEN_273_0; // @[dpath.scala 356:20]
  wire  csr__GEN_456_0; // @[dpath.scala 356:20]
  wire  csr__GEN_351_1; // @[dpath.scala 356:20]
  wire  csr__GEN_450_0; // @[dpath.scala 356:20]
  wire  csr__GEN_357_0; // @[dpath.scala 356:20]
  wire  csr__GEN_279_0; // @[dpath.scala 356:20]
  wire  csr__GEN_399_0; // @[dpath.scala 356:20]
  wire  csr__GEN_264_0; // @[dpath.scala 356:20]
  wire  csr__GEN_300_0; // @[dpath.scala 356:20]
  wire  csr__GEN_432_0; // @[dpath.scala 356:20]
  wire  csr__GEN_381_0; // @[dpath.scala 356:20]
  wire  csr__GEN_339_1; // @[dpath.scala 356:20]
  wire  csr__GEN_261_0; // @[dpath.scala 356:20]
  wire  csr__GEN_360_0; // @[dpath.scala 356:20]
  wire  csr__GEN_246_1; // @[dpath.scala 356:20]
  wire  csr__GEN_438_0; // @[dpath.scala 356:20]
  wire  csr__GEN_282_0; // @[dpath.scala 356:20]
  wire  csr__GEN_345_1; // @[dpath.scala 356:20]
  wire  csr__GEN_240_1; // @[dpath.scala 356:20]
  wire  csr__GEN_444_0; // @[dpath.scala 356:20]
  wire  csr__GEN_267_1; // @[dpath.scala 356:20]
  wire  csr__GEN_459_0; // @[dpath.scala 356:20]
  wire  csr__GEN_453_0; // @[dpath.scala 356:20]
  wire  csr__GEN_366_0; // @[dpath.scala 356:20]
  wire  csr__GEN_7_0; // @[dpath.scala 356:20]
  wire  csr__GEN_324_1; // @[dpath.scala 356:20]
  wire  csr__GEN_333_1; // @[dpath.scala 356:20]
  wire  csr__GEN_342_0; // @[dpath.scala 356:20]
  wire  csr__GEN_405_0; // @[dpath.scala 356:20]
  wire  csr__GEN_420_1; // @[dpath.scala 356:20]
  wire  csr__GEN_306_0; // @[dpath.scala 356:20]
  wire  csr__GEN_3_0; // @[dpath.scala 356:20]
  wire  csr__GEN_426_0; // @[dpath.scala 356:20]
  wire  csr__GEN_441_0; // @[dpath.scala 356:20]
  wire  csr__GEN_348_0; // @[dpath.scala 356:20]
  wire  csr__GEN_255_0; // @[dpath.scala 356:20]
  wire  csr__GEN_146_0; // @[dpath.scala 356:20]
  wire  csr__GEN_363_0; // @[dpath.scala 356:20]
  wire  csr__GEN_321_1; // @[dpath.scala 356:20]
  wire  csr__GEN_327_1; // @[dpath.scala 356:20]
  wire  csr__GEN_354_0; // @[dpath.scala 356:20]
  wire  csr__GEN_234_1; // @[dpath.scala 356:20]
  wire  csr__GEN_249_1; // @[dpath.scala 356:20]
  wire  csr__GEN_243_0; // @[dpath.scala 356:20]
  wire  csr__GEN_447_0; // @[dpath.scala 356:20]
  wire  csr__GEN_330_1; // @[dpath.scala 356:20]
  wire  csr__GEN_429_0; // @[dpath.scala 356:20]
  wire  csr__GEN_293_1; // @[dpath.scala 356:20]
  wire  csr__GEN_414_1; // @[dpath.scala 356:20]
  wire  csr__GEN_309_0; // @[dpath.scala 356:20]
  wire  csr__GEN_299_1; // @[dpath.scala 356:20]
  wire  csr__GEN_336_0; // @[dpath.scala 356:20]
  wire  csr__GEN_408_0; // @[dpath.scala 356:20]
  wire  csr__GEN_150_0; // @[dpath.scala 356:20]
  wire  csr__GEN_435_0; // @[dpath.scala 356:20]
  wire  csr__GEN_392_1; // @[dpath.scala 356:20]
  wire  csr__GEN_398_1; // @[dpath.scala 356:20]
  wire  csr__GEN_423_1; // @[dpath.scala 356:20]
  wire  csr__GEN_237_0; // @[dpath.scala 356:20]
  wire  csr__GEN_315_1; // @[dpath.scala 356:20]
  wire  csr__GEN_302_1; // @[dpath.scala 356:20]
  wire  csr__GEN_380_1; // @[dpath.scala 356:20]
  wire  csr__GEN_318_1; // @[dpath.scala 356:20]
  wire  csr__GEN_287_1; // @[dpath.scala 356:20]
  wire  csr__GEN_386_1; // @[dpath.scala 356:20]
  wire  csr__GEN_281_1; // @[dpath.scala 356:20]
  wire  csr__GEN_312_1; // @[dpath.scala 356:20]
  wire  csr__GEN_417_1; // @[dpath.scala 356:20]
  wire  csr__GEN_411_1; // @[dpath.scala 356:20]
  wire  csr__GEN_401_1; // @[dpath.scala 356:20]
  wire  csr__GEN_374_1; // @[dpath.scala 356:20]
  wire  csr__GEN_368_1; // @[dpath.scala 356:20]
  wire  csr__GEN_383_1; // @[dpath.scala 356:20]
  wire  csr__GEN_263_1; // @[dpath.scala 356:20]
  wire  csr__GEN_446_0; // @[dpath.scala 356:20]
  wire  csr__GEN_290_1; // @[dpath.scala 356:20]
  wire  csr__GEN_389_1; // @[dpath.scala 356:20]
  wire  csr__GEN_254_1; // @[dpath.scala 356:20]
  wire  csr__GEN_461_0; // @[dpath.scala 356:20]
  wire  csr__GEN_362_1; // @[dpath.scala 356:20]
  wire  csr__GEN_296_1; // @[dpath.scala 356:20]
  wire  csr__GEN_395_1; // @[dpath.scala 356:20]
  wire  csr__GEN_275_1; // @[dpath.scala 356:20]
  wire  csr__GEN_269_1; // @[dpath.scala 356:20]
  wire  csr__GEN_278_1; // @[dpath.scala 356:20]
  wire  csr__GEN_251_1; // @[dpath.scala 356:20]
  wire  csr__GEN_455_0; // @[dpath.scala 356:20]
  wire  csr__GEN_377_1; // @[dpath.scala 356:20]
  wire  csr__GEN_272_1; // @[dpath.scala 356:20]
  wire  csr__GEN_335_1; // @[dpath.scala 356:20]
  wire  csr__GEN_434_0; // @[dpath.scala 356:20]
  wire  csr__GEN_257_1; // @[dpath.scala 356:20]
  wire  csr__GEN_443_0; // @[dpath.scala 356:20]
  wire  csr__GEN_356_1; // @[dpath.scala 356:20]
  wire  csr__GEN_350_1; // @[dpath.scala 356:20]
  wire  csr__GEN_428_0; // @[dpath.scala 356:20]
  wire  csr__GEN_449_0; // @[dpath.scala 356:20]
  wire  csr__GEN_236_1; // @[dpath.scala 356:20]
  wire  csr__GEN_371_1; // @[dpath.scala 356:20]
  wire  csr__GEN_284_1; // @[dpath.scala 356:20]
  wire  csr__GEN_416_1; // @[dpath.scala 356:20]
  wire  csr__GEN_260_1; // @[dpath.scala 356:20]
  wire  csr__GEN_338_1; // @[dpath.scala 356:20]
  wire  csr__GEN_344_1; // @[dpath.scala 356:20]
  wire  csr__GEN_239_1; // @[dpath.scala 356:20]
  wire  csr__GEN_353_1; // @[dpath.scala 356:20]
  wire  csr__GEN_266_1; // @[dpath.scala 356:20]
  wire  csr__GEN_452_0; // @[dpath.scala 356:20]
  wire  csr__GEN_365_1; // @[dpath.scala 356:20]
  wire  csr__GEN_6_0; // @[dpath.scala 356:20]
  wire  csr__GEN_410_1; // @[dpath.scala 356:20]
  wire  csr__GEN_152_1; // @[dpath.scala 356:20]
  wire  csr__GEN_437_0; // @[dpath.scala 356:20]
  wire  csr__GEN_332_1; // @[dpath.scala 356:20]
  wire  csr__GEN_245_1; // @[dpath.scala 356:20]
  wire  csr__GEN_359_1; // @[dpath.scala 356:20]
  wire  csr__GEN_431_0; // @[dpath.scala 356:20]
  wire  csr__GEN_458_0; // @[dpath.scala 356:20]
  wire  csr__GEN_317_1; // @[dpath.scala 356:20]
  wire  csr__GEN_326_1; // @[dpath.scala 356:20]
  wire  csr__GEN_341_1; // @[dpath.scala 356:20]
  wire  csr__GEN_394_1; // @[dpath.scala 356:20]
  wire  csr__GEN_248_1; // @[dpath.scala 356:20]
  wire  csr__GEN_347_1; // @[dpath.scala 356:20]
  wire  csr__GEN_425_1; // @[dpath.scala 356:20]
  wire  csr__GEN_305_1; // @[dpath.scala 356:20]
  wire  csr__GEN_419_1; // @[dpath.scala 356:20]
  wire  csr__GEN_320_1; // @[dpath.scala 356:20]
  wire  csr__GEN_413_1; // @[dpath.scala 356:20]
  wire  csr__GEN_440_0; // @[dpath.scala 356:20]
  wire  csr__GEN_295_1; // @[dpath.scala 356:20]
  wire  csr__GEN_404_1; // @[dpath.scala 356:20]
  wire  csr__GEN_403_1; // @[dpath.scala 356:20]
  wire  csr__GEN_242_1; // @[dpath.scala 356:20]
  wire  csr__GEN_15_1; // @[dpath.scala 356:20]
  wire  csr__GEN_308_1; // @[dpath.scala 356:20]
  wire  csr__GEN_149_1; // @[dpath.scala 356:20]
  wire  csr__GEN_329_1; // @[dpath.scala 356:20]
  wire  csr__GEN_292_1; // @[dpath.scala 356:20]
  wire  csr__GEN_298_1; // @[dpath.scala 356:20]
  wire  csr__GEN_391_1; // @[dpath.scala 356:20]
  wire  csr__GEN_314_1; // @[dpath.scala 356:20]
  wire  csr__GEN_323_1; // @[dpath.scala 356:20]
  wire  csr__GEN_376_1; // @[dpath.scala 356:20]
  wire  csr__GEN_422_1; // @[dpath.scala 356:20]
  wire  csr__GEN_277_1; // @[dpath.scala 356:20]
  wire  csr__GEN_407_1; // @[dpath.scala 356:20]
  wire  csr__GEN_397_1; // @[dpath.scala 356:20]
  wire  csr__GEN_379_1; // @[dpath.scala 356:20]
  wire  csr__GEN_373_1; // @[dpath.scala 356:20]
  wire  csr__GEN_364_1; // @[dpath.scala 356:20]
  wire  csr__GEN_259_1; // @[dpath.scala 356:20]
  wire  csr__GEN_265_1; // @[dpath.scala 356:20]
  wire  csr__GEN_301_1; // @[dpath.scala 356:20]
  wire  csr__GEN_286_1; // @[dpath.scala 356:20]
  wire  csr__GEN_400_1; // @[dpath.scala 356:20]
  wire  csr__GEN_358_1; // @[dpath.scala 356:20]
  wire  csr__GEN_385_1; // @[dpath.scala 356:20]
  wire  csr__GEN_457_0; // @[dpath.scala 356:20]
  wire  csr__GEN_311_1; // @[dpath.scala 356:20]
  wire  csr__GEN_280_1; // @[dpath.scala 356:20]
  wire  csr__GEN_367_1; // @[dpath.scala 356:20]
  wire  csr__GEN_247_1; // @[dpath.scala 356:20]
  wire  csr__GEN_274_1; // @[dpath.scala 356:20]
  wire  csr__GEN_460_0; // @[dpath.scala 356:20]
  wire  csr__GEN_283_1; // @[dpath.scala 356:20]
  wire  csr__GEN_388_1; // @[dpath.scala 356:20]
  wire  csr__GEN_382_1; // @[dpath.scala 356:20]
  wire  csr__GEN_268_1; // @[dpath.scala 356:20]
  wire  csr__GEN_346_1; // @[dpath.scala 356:20]
  wire  csr__GEN_340_1; // @[dpath.scala 356:20]
  wire  csr__GEN_439_0; // @[dpath.scala 356:20]
  wire  csr__GEN_262_1; // @[dpath.scala 356:20]
  wire  csr__GEN_361_1; // @[dpath.scala 356:20]
  wire  csr__GEN_241_1; // @[dpath.scala 356:20]
  wire  csr__GEN_445_0; // @[dpath.scala 356:20]
  wire  csr__GEN_289_1; // @[dpath.scala 356:20]
  wire  csr__GEN_421_1; // @[dpath.scala 356:20]
  wire  csr__GEN_427_0; // @[dpath.scala 356:20]
  wire  csr__GEN_454_0; // @[dpath.scala 356:20]
  wire  csr__GEN_256_1; // @[dpath.scala 356:20]
  wire  csr__GEN_5_2; // @[dpath.scala 356:20]
  wire  csr__GEN_271_1; // @[dpath.scala 356:20]
  wire  csr__GEN_322_1; // @[dpath.scala 356:20]
  wire  csr__GEN_334_1; // @[dpath.scala 356:20]
  wire  csr__GEN_235_1; // @[dpath.scala 356:20]
  wire  csr__GEN_349_1; // @[dpath.scala 356:20]
  wire  csr__GEN_147_2; // @[dpath.scala 356:20]
  wire  csr__GEN_448_0; // @[dpath.scala 356:20]
  wire  csr__GEN_442_0; // @[dpath.scala 356:20]
  wire  csr__GEN_343_1; // @[dpath.scala 356:20]
  wire  csr__GEN_355_1; // @[dpath.scala 356:20]
  wire  csr__GEN_370_1; // @[dpath.scala 356:20]
  wire  csr__GEN_250_1; // @[dpath.scala 356:20]
  wire  csr__GEN_463_0; // @[dpath.scala 356:20]
  wire  csr__GEN_328_1; // @[dpath.scala 356:20]
  reg [31:0] if_reg_pc; // @[dpath.scala 52:35]
  reg [31:0] dec_reg_inst; // @[dpath.scala 55:35]
  reg [31:0] dec_reg_pc; // @[dpath.scala 56:35]
  reg [31:0] exe_reg_inst; // @[dpath.scala 59:35]
  reg [31:0] exe_reg_pc; // @[dpath.scala 60:35]
  reg [4:0] exe_reg_wbaddr; // @[dpath.scala 61:35]
  reg [31:0] exe_alu_op1; // @[dpath.scala 64:35]
  reg [31:0] brjmp_offset; // @[dpath.scala 65:35]
  reg [31:0] exe_reg_rs2_data; // @[dpath.scala 66:35]
  reg [3:0] exe_reg_ctrl_br_type; // @[dpath.scala 67:35]
  reg [3:0] exe_reg_ctrl_alu_fun; // @[dpath.scala 69:35]
  reg [1:0] exe_reg_ctrl_wb_sel; // @[dpath.scala 70:35]
  reg  exe_reg_ctrl_rf_wen; // @[dpath.scala 71:35]
  reg  exe_reg_ctrl_mem_val; // @[dpath.scala 72:35]
  reg  exe_reg_ctrl_mem_fcn; // @[dpath.scala 73:35]
  reg [2:0] exe_reg_ctrl_mem_typ; // @[dpath.scala 74:35]
  reg [2:0] exe_reg_ctrl_csr_cmd; // @[dpath.scala 75:35]
  reg [31:0] mem_reg_pc; // @[dpath.scala 78:35]
  reg [31:0] mem_reg_inst; // @[dpath.scala 79:35]
  reg [31:0] mem_reg_alu_out; // @[dpath.scala 80:35]
  reg [4:0] mem_reg_wbaddr; // @[dpath.scala 81:35]
  reg [31:0] mem_reg_rs2_data; // @[dpath.scala 86:35]
  reg  mem_reg_ctrl_rf_wen; // @[dpath.scala 87:35]
  reg  mem_reg_ctrl_mem_val; // @[dpath.scala 88:35]
  reg  mem_reg_ctrl_mem_fcn; // @[dpath.scala 89:35]
  reg [2:0] mem_reg_ctrl_mem_typ; // @[dpath.scala 90:35]
  reg [1:0] mem_reg_ctrl_wb_sel; // @[dpath.scala 91:35]
  reg [2:0] mem_reg_ctrl_csr_cmd; // @[dpath.scala 92:35]
  reg [4:0] wb_reg_wbaddr; // @[dpath.scala 95:35]
  reg [31:0] wb_reg_wbdata; // @[dpath.scala 96:35]
  reg  wb_reg_ctrl_rf_wen; // @[dpath.scala 97:35]
  wire  _T_145 = ~io_ctl_dec_stall; // @[dpath.scala 107:11]
  wire  _T_147 = ~io_ctl_full_stall; // @[dpath.scala 107:32]
  wire  _T_148 = _T_145 & _T_147; // @[dpath.scala 107:29]
  wire  _T_149 = _T_148 | io_ctl_pipeline_kill; // @[dpath.scala 107:52]
  wire  _T_158 = io_ctl_exe_pc_sel == 2'h0; // @[dpath.scala 120:45]
  wire  _T_159 = io_ctl_fencei & _T_158; // @[dpath.scala 120:24]
  wire  _T_162 = _T_159 & _T_145; // @[dpath.scala 120:54]
  wire  _T_165 = _T_162 & _T_147; // @[dpath.scala 121:28]
  wire  _T_167 = ~io_ctl_pipeline_kill; // @[dpath.scala 121:53]
  wire  _T_168 = _T_165 & _T_167; // @[dpath.scala 121:50]
  wire [31:0] if_pc_plus4 = if_reg_pc + 32'h4; // @[dpath.scala 112:33]
  wire  _T_153 = io_ctl_exe_pc_sel == 2'h1; // @[dpath.scala 115:40]
  wire [31:0] exe_brjmp_target = exe_reg_pc + brjmp_offset; // @[dpath.scala 320:38]
  wire  _T_154 = io_ctl_exe_pc_sel == 2'h2; // @[dpath.scala 116:40]
  wire [31:0] exe_adder_out = exe_alu_op1 + brjmp_offset; // @[dpath.scala 300:37]
  wire [31:0] exception_target = csr_io_evec; // @[dpath.scala 105:34 dpath.scala 365:21]
  wire [4:0] dec_rs1_addr = dec_reg_inst[19:15]; // @[dpath.scala 151:35]
  wire [4:0] dec_rs2_addr = dec_reg_inst[24:20]; // @[dpath.scala 152:35]
  wire [4:0] dec_wbaddr = dec_reg_inst[11:7]; // @[dpath.scala 153:35]
  wire [11:0] imm_itype = dec_reg_inst[31:20]; // @[dpath.scala 174:33]
  wire [11:0] imm_stype = {dec_reg_inst[31:25],dec_wbaddr}; // @[Cat.scala 30:58]
  wire [11:0] imm_sbtype = {dec_reg_inst[31],dec_reg_inst[7],dec_reg_inst[30:25],dec_reg_inst[11:8]}; // @[Cat.scala 30:58]
  wire [19:0] imm_utype = dec_reg_inst[31:12]; // @[dpath.scala 177:33]
  wire [19:0] imm_ujtype = {dec_reg_inst[31],dec_reg_inst[19:12],dec_reg_inst[20],dec_reg_inst[30:21]}; // @[Cat.scala 30:58]
  wire [31:0] imm_z = {27'h0,dec_rs1_addr}; // @[Cat.scala 30:58]
  wire [19:0] _T_198 = imm_itype[11] ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire [31:0] imm_itype_sext = {_T_198,imm_itype}; // @[Cat.scala 30:58]
  wire [19:0] _T_203 = imm_stype[11] ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire [31:0] imm_stype_sext = {_T_203,dec_reg_inst[31:25],dec_wbaddr}; // @[Cat.scala 30:58]
  wire [18:0] _T_208 = imm_sbtype[11] ? 19'h7ffff : 19'h0; // @[Bitwise.scala 72:12]
  wire [31:0] imm_sbtype_sext = {_T_208,dec_reg_inst[31],dec_reg_inst[7],dec_reg_inst[30:25],dec_reg_inst[11:8],1'h0}; // @[Cat.scala 30:58]
  wire [31:0] imm_utype_sext = {imm_utype,12'h0}; // @[Cat.scala 30:58]
  wire [10:0] _T_220 = imm_ujtype[19] ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [31:0] imm_ujtype_sext = {_T_220,dec_reg_inst[31],dec_reg_inst[19:12],dec_reg_inst[20],dec_reg_inst[30:21],1'h0}; // @[Cat.scala 30:58]
  wire  _T_224 = io_ctl_op2_sel == 3'h0; // @[dpath.scala 191:32]
  wire  _T_225 = io_ctl_op2_sel == 3'h1; // @[dpath.scala 192:32]
  wire  _T_226 = io_ctl_op2_sel == 3'h2; // @[dpath.scala 193:32]
  wire  _T_227 = io_ctl_op2_sel == 3'h3; // @[dpath.scala 194:32]
  wire  _T_228 = io_ctl_op2_sel == 3'h4; // @[dpath.scala 195:32]
  wire  _T_229 = io_ctl_op2_sel == 3'h5; // @[dpath.scala 196:32]
  wire  _T_240 = io_ctl_op1_sel == 2'h2; // @[dpath.scala 213:45]
  wire  _T_241 = io_ctl_op1_sel == 2'h1; // @[dpath.scala 214:45]
  wire  _T_242 = exe_reg_wbaddr == dec_rs1_addr; // @[dpath.scala 215:45]
  wire  _T_244 = dec_rs1_addr != 5'h0; // @[dpath.scala 215:80]
  wire  _T_245 = _T_242 & _T_244; // @[dpath.scala 215:63]
  wire  _T_246 = _T_245 & exe_reg_ctrl_rf_wen; // @[dpath.scala 215:88]
  wire  _T_247 = mem_reg_wbaddr == dec_rs1_addr; // @[dpath.scala 216:45]
  wire  _T_250 = _T_247 & _T_244; // @[dpath.scala 216:63]
  wire  _T_251 = _T_250 & mem_reg_ctrl_rf_wen; // @[dpath.scala 216:88]
  wire  _T_252 = wb_reg_wbaddr == dec_rs1_addr; // @[dpath.scala 217:45]
  wire  _T_255 = _T_252 & _T_244; // @[dpath.scala 217:63]
  wire  _T_256 = _T_255 & wb_reg_ctrl_rf_wen; // @[dpath.scala 217:88]
  wire  _T_439 = mem_reg_ctrl_wb_sel == 2'h0; // @[dpath.scala 376:40]
  wire  _T_440 = mem_reg_ctrl_wb_sel == 2'h2; // @[dpath.scala 377:40]
  wire  _T_441 = mem_reg_ctrl_wb_sel == 2'h1; // @[dpath.scala 378:40]
  wire  _T_442 = mem_reg_ctrl_wb_sel == 2'h3; // @[dpath.scala 379:40]
  wire  _T_321 = exe_reg_ctrl_alu_fun == 4'h0; // @[dpath.scala 304:41]
  wire  _T_322 = exe_reg_ctrl_alu_fun == 4'h1; // @[dpath.scala 305:41]
  wire [31:0] _T_325 = exe_alu_op1 - brjmp_offset; // @[dpath.scala 305:71]
  wire  _T_326 = exe_reg_ctrl_alu_fun == 4'h5; // @[dpath.scala 306:41]
  wire [31:0] _T_327 = exe_alu_op1 & brjmp_offset; // @[dpath.scala 306:71]
  wire  _T_328 = exe_reg_ctrl_alu_fun == 4'h6; // @[dpath.scala 307:41]
  wire [31:0] _T_329 = exe_alu_op1 | brjmp_offset; // @[dpath.scala 307:71]
  wire  _T_330 = exe_reg_ctrl_alu_fun == 4'h7; // @[dpath.scala 308:41]
  wire [31:0] _T_331 = exe_alu_op1 ^ brjmp_offset; // @[dpath.scala 308:71]
  wire  _T_332 = exe_reg_ctrl_alu_fun == 4'h8; // @[dpath.scala 309:41]
  wire  _T_335 = $signed(exe_alu_op1) < $signed(brjmp_offset); // @[dpath.scala 309:78]
  wire  _T_336 = exe_reg_ctrl_alu_fun == 4'h9; // @[dpath.scala 310:41]
  wire  _T_337 = exe_alu_op1 < brjmp_offset; // @[dpath.scala 310:71]
  wire  _T_338 = exe_reg_ctrl_alu_fun == 4'h2; // @[dpath.scala 311:41]
  wire [4:0] alu_shamt = brjmp_offset[4:0]; // @[dpath.scala 299:35]
  wire [62:0] _GEN_84 = {{31'd0}, exe_alu_op1}; // @[dpath.scala 311:72]
  wire [62:0] _T_339 = _GEN_84 << alu_shamt; // @[dpath.scala 311:72]
  wire  _T_341 = exe_reg_ctrl_alu_fun == 4'h4; // @[dpath.scala 312:41]
  wire [31:0] _T_344 = $signed(exe_alu_op1) >>> alu_shamt;
  wire  _T_345 = exe_reg_ctrl_alu_fun == 4'h3; // @[dpath.scala 313:41]
  wire [31:0] _T_346 = exe_alu_op1 >> alu_shamt; // @[dpath.scala 313:71]
  wire  _T_347 = exe_reg_ctrl_alu_fun == 4'ha; // @[dpath.scala 314:41]
  wire  _T_348 = exe_reg_ctrl_alu_fun == 4'hb; // @[dpath.scala 315:41]
  wire  _T_262 = exe_reg_wbaddr == dec_rs2_addr; // @[dpath.scala 221:45]
  wire  _T_264 = dec_rs2_addr != 5'h0; // @[dpath.scala 221:80]
  wire  _T_265 = _T_262 & _T_264; // @[dpath.scala 221:63]
  wire  _T_266 = _T_265 & exe_reg_ctrl_rf_wen; // @[dpath.scala 221:88]
  wire  _T_268 = _T_266 & _T_224; // @[dpath.scala 221:111]
  wire  _T_269 = mem_reg_wbaddr == dec_rs2_addr; // @[dpath.scala 222:45]
  wire  _T_272 = _T_269 & _T_264; // @[dpath.scala 222:63]
  wire  _T_273 = _T_272 & mem_reg_ctrl_rf_wen; // @[dpath.scala 222:88]
  wire  _T_275 = _T_273 & _T_224; // @[dpath.scala 222:111]
  wire  _T_276 = wb_reg_wbaddr == dec_rs2_addr; // @[dpath.scala 223:45]
  wire  _T_279 = _T_276 & _T_264; // @[dpath.scala 223:63]
  wire  _T_280 = _T_279 & wb_reg_ctrl_rf_wen; // @[dpath.scala 223:88]
  wire  _T_282 = _T_280 & _T_224; // @[dpath.scala 223:111]
  wire  _T_306 = io_ctl_dec_stall & _T_147; // @[dpath.scala 244:28]
  wire  _T_307 = _T_306 | io_ctl_pipeline_kill; // @[dpath.scala 244:51]
  wire [1:0] _GEN_11 = io_ctl_dec_kill ? 2'h0 : io_ctl_mem_fcn; // @[dpath.scala 270:7]
  wire [1:0] _GEN_28 = _T_148 ? _GEN_11 : {{1'd0}, exe_reg_ctrl_mem_fcn}; // @[dpath.scala 257:4]
  wire [1:0] _GEN_36 = _T_307 ? 2'h0 : _GEN_28; // @[dpath.scala 245:4]
  wire [31:0] exe_pc_plus4 = exe_reg_pc + 32'h4; // @[dpath.scala 323:38]
  wire  _T_371 = exe_reg_ctrl_wb_sel == 2'h2; // @[dpath.scala 336:57]
  wire  _T_450 = io_ctl_mem_exception ? 1'h0 : mem_reg_ctrl_rf_wen; // @[dpath.scala 390:34]
  wire  _GEN_81 = _T_147 & _T_450; // @[dpath.scala 387:4]
  RegisterFile regfile ( // @[dpath.scala 157:24]
    .metaReset(regfile_metaReset),
    .clock(regfile_clock),
    .io_rs1_addr(regfile_io_rs1_addr),
    .io_rs1_data(regfile_io_rs1_data),
    .io_rs2_addr(regfile_io_rs2_addr),
    .io_rs2_data(regfile_io_rs2_data),
    .io_waddr(regfile_io_waddr),
    .io_wdata(regfile_io_wdata),
    .io_wen(regfile_io_wen),
    ._GEN_0_0(regfile__GEN_0_0),
    ._GEN_1_3(regfile__GEN_1_3)
  );
  CSRFile csr ( // @[dpath.scala 356:20]
    .metaReset(csr_metaReset),
    .clock(csr_clock),
    .reset(csr_reset),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_eret(csr_io_eret),
    .io_decode_csr(csr_io_decode_csr),
    .io_status_debug(csr_io_status_debug),
    .io_status_prv(csr_io_status_prv),
    .io_status_sd(csr_io_status_sd),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_tsr(csr_io_status_tsr),
    .io_status_tw(csr_io_status_tw),
    .io_status_tvm(csr_io_status_tvm),
    .io_status_mxr(csr_io_status_mxr),
    .io_status_sum(csr_io_status_sum),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_xs(csr_io_status_xs),
    .io_status_fs(csr_io_status_fs),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_hpp(csr_io_status_hpp),
    .io_status_spp(csr_io_status_spp),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_hpie(csr_io_status_hpie),
    .io_status_spie(csr_io_status_spie),
    .io_status_upie(csr_io_status_upie),
    .io_status_mie(csr_io_status_mie),
    .io_status_hie(csr_io_status_hie),
    .io_status_sie(csr_io_status_sie),
    .io_status_uie(csr_io_status_uie),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_retire(csr_io_retire),
    .io_pc(csr_io_pc),
    ._GEN_451_0(csr__GEN_451_0),
    ._GEN_331_0(csr__GEN_331_0),
    ._GEN_337_0(csr__GEN_337_0),
    ._GEN_415_0(csr__GEN_415_0),
    ._GEN_436_0(csr__GEN_436_0),
    ._GEN_352_0(csr__GEN_352_0),
    ._GEN_430_0(csr__GEN_430_0),
    ._GEN_151_0(csr__GEN_151_0),
    ._GEN_310_0(csr__GEN_310_0),
    ._GEN_409_0(csr__GEN_409_0),
    ._GEN_253_0(csr__GEN_253_0),
    ._GEN_316_0(csr__GEN_316_0),
    ._GEN_244_0(csr__GEN_244_0),
    ._GEN_238_0(csr__GEN_238_0),
    ._GEN_325_0(csr__GEN_325_0),
    ._GEN_433_0(csr__GEN_433_0),
    ._GEN_313_0(csr__GEN_313_0),
    ._GEN_11_0(csr__GEN_11_0),
    ._GEN_304_0(csr__GEN_304_0),
    ._GEN_294_0(csr__GEN_294_0),
    ._GEN_303_0(csr__GEN_303_0),
    ._GEN_402_0(csr__GEN_402_0),
    ._GEN_412_0(csr__GEN_412_0),
    ._GEN_424_0(csr__GEN_424_0),
    ._GEN_319_0(csr__GEN_319_0),
    ._GEN_288_0(csr__GEN_288_0),
    ._GEN_418_0(csr__GEN_418_0),
    ._GEN_387_0(csr__GEN_387_0),
    ._GEN_462_0(csr__GEN_462_0),
    ._GEN_375_0(csr__GEN_375_0),
    ._GEN_390_0(csr__GEN_390_0),
    ._GEN_307_0(csr__GEN_307_0),
    ._GEN_297_0(csr__GEN_297_0),
    ._GEN_406_0(csr__GEN_406_0),
    ._GEN_270_0(csr__GEN_270_0),
    ._GEN_369_0(csr__GEN_369_0),
    ._GEN_396_0(csr__GEN_396_0),
    ._GEN_276_0(csr__GEN_276_0),
    ._GEN_291_0(csr__GEN_291_0),
    ._GEN_258_0(csr__GEN_258_0),
    ._GEN_372_0(csr__GEN_372_0),
    ._GEN_252_1(csr__GEN_252_1),
    ._GEN_285_0(csr__GEN_285_0),
    ._GEN_384_0(csr__GEN_384_0),
    ._GEN_378_0(csr__GEN_378_0),
    ._GEN_393_0(csr__GEN_393_0),
    ._GEN_273_0(csr__GEN_273_0),
    ._GEN_456_0(csr__GEN_456_0),
    ._GEN_351_1(csr__GEN_351_1),
    ._GEN_450_0(csr__GEN_450_0),
    ._GEN_357_0(csr__GEN_357_0),
    ._GEN_279_0(csr__GEN_279_0),
    ._GEN_399_0(csr__GEN_399_0),
    ._GEN_264_0(csr__GEN_264_0),
    ._GEN_300_0(csr__GEN_300_0),
    ._GEN_432_0(csr__GEN_432_0),
    ._GEN_381_0(csr__GEN_381_0),
    ._GEN_339_1(csr__GEN_339_1),
    ._GEN_261_0(csr__GEN_261_0),
    ._GEN_360_0(csr__GEN_360_0),
    ._GEN_246_1(csr__GEN_246_1),
    ._GEN_438_0(csr__GEN_438_0),
    ._GEN_282_0(csr__GEN_282_0),
    ._GEN_345_1(csr__GEN_345_1),
    ._GEN_240_1(csr__GEN_240_1),
    ._GEN_444_0(csr__GEN_444_0),
    ._GEN_267_1(csr__GEN_267_1),
    ._GEN_459_0(csr__GEN_459_0),
    ._GEN_453_0(csr__GEN_453_0),
    ._GEN_366_0(csr__GEN_366_0),
    ._GEN_7_0(csr__GEN_7_0),
    ._GEN_324_1(csr__GEN_324_1),
    ._GEN_333_1(csr__GEN_333_1),
    ._GEN_342_0(csr__GEN_342_0),
    ._GEN_405_0(csr__GEN_405_0),
    ._GEN_420_1(csr__GEN_420_1),
    ._GEN_306_0(csr__GEN_306_0),
    ._GEN_3_0(csr__GEN_3_0),
    ._GEN_426_0(csr__GEN_426_0),
    ._GEN_441_0(csr__GEN_441_0),
    ._GEN_348_0(csr__GEN_348_0),
    ._GEN_255_0(csr__GEN_255_0),
    ._GEN_146_0(csr__GEN_146_0),
    ._GEN_363_0(csr__GEN_363_0),
    ._GEN_321_1(csr__GEN_321_1),
    ._GEN_327_1(csr__GEN_327_1),
    ._GEN_354_0(csr__GEN_354_0),
    ._GEN_234_1(csr__GEN_234_1),
    ._GEN_249_1(csr__GEN_249_1),
    ._GEN_243_0(csr__GEN_243_0),
    ._GEN_447_0(csr__GEN_447_0),
    ._GEN_330_1(csr__GEN_330_1),
    ._GEN_429_0(csr__GEN_429_0),
    ._GEN_293_1(csr__GEN_293_1),
    ._GEN_414_1(csr__GEN_414_1),
    ._GEN_309_0(csr__GEN_309_0),
    ._GEN_299_1(csr__GEN_299_1),
    ._GEN_336_0(csr__GEN_336_0),
    ._GEN_408_0(csr__GEN_408_0),
    ._GEN_150_0(csr__GEN_150_0),
    ._GEN_435_0(csr__GEN_435_0),
    ._GEN_392_1(csr__GEN_392_1),
    ._GEN_398_1(csr__GEN_398_1),
    ._GEN_423_1(csr__GEN_423_1),
    ._GEN_237_0(csr__GEN_237_0),
    ._GEN_315_1(csr__GEN_315_1),
    ._GEN_302_1(csr__GEN_302_1),
    ._GEN_380_1(csr__GEN_380_1),
    ._GEN_318_1(csr__GEN_318_1),
    ._GEN_287_1(csr__GEN_287_1),
    ._GEN_386_1(csr__GEN_386_1),
    ._GEN_281_1(csr__GEN_281_1),
    ._GEN_312_1(csr__GEN_312_1),
    ._GEN_417_1(csr__GEN_417_1),
    ._GEN_411_1(csr__GEN_411_1),
    ._GEN_401_1(csr__GEN_401_1),
    ._GEN_374_1(csr__GEN_374_1),
    ._GEN_368_1(csr__GEN_368_1),
    ._GEN_383_1(csr__GEN_383_1),
    ._GEN_263_1(csr__GEN_263_1),
    ._GEN_446_0(csr__GEN_446_0),
    ._GEN_290_1(csr__GEN_290_1),
    ._GEN_389_1(csr__GEN_389_1),
    ._GEN_254_1(csr__GEN_254_1),
    ._GEN_461_0(csr__GEN_461_0),
    ._GEN_362_1(csr__GEN_362_1),
    ._GEN_296_1(csr__GEN_296_1),
    ._GEN_395_1(csr__GEN_395_1),
    ._GEN_275_1(csr__GEN_275_1),
    ._GEN_269_1(csr__GEN_269_1),
    ._GEN_278_1(csr__GEN_278_1),
    ._GEN_251_1(csr__GEN_251_1),
    ._GEN_455_0(csr__GEN_455_0),
    ._GEN_377_1(csr__GEN_377_1),
    ._GEN_272_1(csr__GEN_272_1),
    ._GEN_335_1(csr__GEN_335_1),
    ._GEN_434_0(csr__GEN_434_0),
    ._GEN_257_1(csr__GEN_257_1),
    ._GEN_443_0(csr__GEN_443_0),
    ._GEN_356_1(csr__GEN_356_1),
    ._GEN_350_1(csr__GEN_350_1),
    ._GEN_428_0(csr__GEN_428_0),
    ._GEN_449_0(csr__GEN_449_0),
    ._GEN_236_1(csr__GEN_236_1),
    ._GEN_371_1(csr__GEN_371_1),
    ._GEN_284_1(csr__GEN_284_1),
    ._GEN_416_1(csr__GEN_416_1),
    ._GEN_260_1(csr__GEN_260_1),
    ._GEN_338_1(csr__GEN_338_1),
    ._GEN_344_1(csr__GEN_344_1),
    ._GEN_239_1(csr__GEN_239_1),
    ._GEN_353_1(csr__GEN_353_1),
    ._GEN_266_1(csr__GEN_266_1),
    ._GEN_452_0(csr__GEN_452_0),
    ._GEN_365_1(csr__GEN_365_1),
    ._GEN_6_0(csr__GEN_6_0),
    ._GEN_410_1(csr__GEN_410_1),
    ._GEN_152_1(csr__GEN_152_1),
    ._GEN_437_0(csr__GEN_437_0),
    ._GEN_332_1(csr__GEN_332_1),
    ._GEN_245_1(csr__GEN_245_1),
    ._GEN_359_1(csr__GEN_359_1),
    ._GEN_431_0(csr__GEN_431_0),
    ._GEN_458_0(csr__GEN_458_0),
    ._GEN_317_1(csr__GEN_317_1),
    ._GEN_326_1(csr__GEN_326_1),
    ._GEN_341_1(csr__GEN_341_1),
    ._GEN_394_1(csr__GEN_394_1),
    ._GEN_248_1(csr__GEN_248_1),
    ._GEN_347_1(csr__GEN_347_1),
    ._GEN_425_1(csr__GEN_425_1),
    ._GEN_305_1(csr__GEN_305_1),
    ._GEN_419_1(csr__GEN_419_1),
    ._GEN_320_1(csr__GEN_320_1),
    ._GEN_413_1(csr__GEN_413_1),
    ._GEN_440_0(csr__GEN_440_0),
    ._GEN_295_1(csr__GEN_295_1),
    ._GEN_404_1(csr__GEN_404_1),
    ._GEN_403_1(csr__GEN_403_1),
    ._GEN_242_1(csr__GEN_242_1),
    ._GEN_15_1(csr__GEN_15_1),
    ._GEN_308_1(csr__GEN_308_1),
    ._GEN_149_1(csr__GEN_149_1),
    ._GEN_329_1(csr__GEN_329_1),
    ._GEN_292_1(csr__GEN_292_1),
    ._GEN_298_1(csr__GEN_298_1),
    ._GEN_391_1(csr__GEN_391_1),
    ._GEN_314_1(csr__GEN_314_1),
    ._GEN_323_1(csr__GEN_323_1),
    ._GEN_376_1(csr__GEN_376_1),
    ._GEN_422_1(csr__GEN_422_1),
    ._GEN_277_1(csr__GEN_277_1),
    ._GEN_407_1(csr__GEN_407_1),
    ._GEN_397_1(csr__GEN_397_1),
    ._GEN_379_1(csr__GEN_379_1),
    ._GEN_373_1(csr__GEN_373_1),
    ._GEN_364_1(csr__GEN_364_1),
    ._GEN_259_1(csr__GEN_259_1),
    ._GEN_265_1(csr__GEN_265_1),
    ._GEN_301_1(csr__GEN_301_1),
    ._GEN_286_1(csr__GEN_286_1),
    ._GEN_400_1(csr__GEN_400_1),
    ._GEN_358_1(csr__GEN_358_1),
    ._GEN_385_1(csr__GEN_385_1),
    ._GEN_457_0(csr__GEN_457_0),
    ._GEN_311_1(csr__GEN_311_1),
    ._GEN_280_1(csr__GEN_280_1),
    ._GEN_367_1(csr__GEN_367_1),
    ._GEN_247_1(csr__GEN_247_1),
    ._GEN_274_1(csr__GEN_274_1),
    ._GEN_460_0(csr__GEN_460_0),
    ._GEN_283_1(csr__GEN_283_1),
    ._GEN_388_1(csr__GEN_388_1),
    ._GEN_382_1(csr__GEN_382_1),
    ._GEN_268_1(csr__GEN_268_1),
    ._GEN_346_1(csr__GEN_346_1),
    ._GEN_340_1(csr__GEN_340_1),
    ._GEN_439_0(csr__GEN_439_0),
    ._GEN_262_1(csr__GEN_262_1),
    ._GEN_361_1(csr__GEN_361_1),
    ._GEN_241_1(csr__GEN_241_1),
    ._GEN_445_0(csr__GEN_445_0),
    ._GEN_289_1(csr__GEN_289_1),
    ._GEN_421_1(csr__GEN_421_1),
    ._GEN_427_0(csr__GEN_427_0),
    ._GEN_454_0(csr__GEN_454_0),
    ._GEN_256_1(csr__GEN_256_1),
    ._GEN_5_2(csr__GEN_5_2),
    ._GEN_271_1(csr__GEN_271_1),
    ._GEN_322_1(csr__GEN_322_1),
    ._GEN_334_1(csr__GEN_334_1),
    ._GEN_235_1(csr__GEN_235_1),
    ._GEN_349_1(csr__GEN_349_1),
    ._GEN_147_2(csr__GEN_147_2),
    ._GEN_448_0(csr__GEN_448_0),
    ._GEN_442_0(csr__GEN_442_0),
    ._GEN_343_1(csr__GEN_343_1),
    ._GEN_355_1(csr__GEN_355_1),
    ._GEN_370_1(csr__GEN_370_1),
    ._GEN_250_1(csr__GEN_250_1),
    ._GEN_463_0(csr__GEN_463_0),
    ._GEN_328_1(csr__GEN_328_1)
  );
  assign regfile_metaReset = metaReset;
  assign csr_metaReset = metaReset;
  assign io_imem_req_bits_addr = if_reg_pc; // @[dpath.scala 127:26]
  assign io_dmem_req_valid = mem_reg_ctrl_mem_val; // @[dpath.scala 412:26]
  assign io_dmem_req_bits_addr = mem_reg_alu_out; // @[dpath.scala 413:26]
  assign io_dmem_req_bits_data = mem_reg_rs2_data; // @[dpath.scala 416:26]
  assign io_dmem_req_bits_fcn = mem_reg_ctrl_mem_fcn; // @[dpath.scala 414:26]
  assign io_dmem_req_bits_typ = mem_reg_ctrl_mem_typ; // @[dpath.scala 415:26]
  assign io_dat_dec_inst = dec_reg_inst; // @[dpath.scala 403:22]
  assign io_dat_exe_br_eq = exe_alu_op1 == exe_reg_rs2_data; // @[dpath.scala 404:22]
  assign io_dat_exe_br_lt = $signed(exe_alu_op1) < $signed(exe_reg_rs2_data); // @[dpath.scala 405:22]
  assign io_dat_exe_br_ltu = exe_alu_op1 < exe_reg_rs2_data; // @[dpath.scala 406:22]
  assign io_dat_exe_br_type = exe_reg_ctrl_br_type; // @[dpath.scala 407:22]
  assign io_dat_mem_ctrl_dmem_val = mem_reg_ctrl_mem_val; // @[dpath.scala 409:29]
  assign io_dat_csr_eret = csr_io_eret; // @[dpath.scala 367:20]
  assign _GEN_451 = csr__GEN_451_0;
  assign _GEN_331 = csr__GEN_331_0;
  assign _GEN_337 = csr__GEN_337_0;
  assign _GEN_113_0 = _T_145 & _T_147;
  assign _GEN_415 = csr__GEN_415_0;
  assign _GEN_436 = csr__GEN_436_0;
  assign _GEN_140_0 = ~io_ctl_full_stall;
  assign _GEN_98_0 = _T_279 & wb_reg_ctrl_rf_wen;
  assign _GEN_352 = csr__GEN_352_0;
  assign _GEN_125_0 = _T_306 | io_ctl_pipeline_kill;
  assign _GEN_430 = csr__GEN_430_0;
  assign _GEN_119_0 = _T_145 & _T_147;
  assign _GEN_88_0 = exe_reg_ctrl_alu_fun == 4'h6;
  assign _GEN_151_0 = csr__GEN_151_0;
  assign _GEN_310 = csr__GEN_310_0;
  assign _GEN_104_0 = io_ctl_dec_kill;
  assign _GEN_409 = csr__GEN_409_0;
  assign _GEN_253 = csr__GEN_253_0;
  assign _GEN_316 = csr__GEN_316_0;
  assign _GEN_244 = csr__GEN_244_0;
  assign _GEN_238 = csr__GEN_238_0;
  assign _GEN_101_0 = io_ctl_dec_kill;
  assign _GEN_325 = csr__GEN_325_0;
  assign _GEN_169_0 = io_ctl_pipeline_kill;
  assign _GEN_433 = csr__GEN_433_0;
  assign _GEN_313 = csr__GEN_313_0;
  assign _GEN_91_0 = exe_reg_ctrl_alu_fun == 4'h0;
  assign _GEN_11_0 = csr__GEN_11_0;
  assign _GEN_304 = csr__GEN_304_0;
  assign _GEN_294 = csr__GEN_294_0;
  assign _GEN_303 = csr__GEN_303_0;
  assign _GEN_107_0 = io_ctl_dec_kill;
  assign _GEN_0_0 = regfile__GEN_0_0;
  assign _GEN_402 = csr__GEN_402_0;
  assign _GEN_412 = csr__GEN_412_0;
  assign _GEN_424 = csr__GEN_424_0;
  assign _GEN_175_0 = io_ctl_pipeline_kill;
  assign _GEN_319 = csr__GEN_319_0;
  assign _GEN_288 = csr__GEN_288_0;
  assign _GEN_56_0 = io_ctl_op2_sel == 3'h3;
  assign _GEN_418 = csr__GEN_418_0;
  assign _GEN_122_0 = _T_145 & _T_147;
  assign _GEN_387 = csr__GEN_387_0;
  assign _GEN_72_0 = mem_reg_ctrl_wb_sel == 2'h1;
  assign _GEN_75_0 = _T_250 & mem_reg_ctrl_rf_wen;
  assign _GEN_85_0 = exe_reg_ctrl_alu_fun == 4'h9;
  assign _GEN_178_0 = ~io_ctl_full_stall;
  assign _GEN_157_0 = _T_306 | io_ctl_pipeline_kill;
  assign _GEN_462 = csr__GEN_462_0;
  assign _GEN_69_0 = io_ctl_op2_sel == 3'h0;
  assign _GEN_375 = csr__GEN_375_0;
  assign _GEN_151_1 = reset;
  assign _GEN_33_0 = _T_148 | io_ctl_pipeline_kill;
  assign _GEN_390 = csr__GEN_390_0;
  assign _GEN_307 = csr__GEN_307_0;
  assign _GEN_297 = csr__GEN_297_0;
  assign _GEN_406 = csr__GEN_406_0;
  assign _GEN_270 = csr__GEN_270_0;
  assign _GEN_95_0 = _T_280 & _T_224;
  assign _GEN_45_0 = imm_itype[11];
  assign _GEN_369 = csr__GEN_369_0;
  assign _GEN_396 = csr__GEN_396_0;
  assign _GEN_172_0 = reset;
  assign _GEN_276 = csr__GEN_276_0;
  assign _GEN_291 = csr__GEN_291_0;
  assign _GEN_258 = csr__GEN_258_0;
  assign _GEN_372 = csr__GEN_372_0;
  assign _GEN_252_0 = csr__GEN_252_1;
  assign _GEN_166_0 = io_ctl_pipeline_kill;
  assign _GEN_285 = csr__GEN_285_0;
  assign _GEN_42_0 = _T_145 & _T_147;
  assign _GEN_384 = csr__GEN_384_0;
  assign _GEN_378 = csr__GEN_378_0;
  assign _GEN_393 = csr__GEN_393_0;
  assign _GEN_273 = csr__GEN_273_0;
  assign _GEN_456 = csr__GEN_456_0;
  assign _GEN_80_0 = exe_reg_ctrl_alu_fun == 4'h3;
  assign _GEN_351_0 = csr__GEN_351_1;
  assign _GEN_139_0 = ~io_ctl_full_stall;
  assign _GEN_145_0 = io_ctl_pipeline_kill;
  assign _GEN_450 = csr__GEN_450_0;
  assign _GEN_53_1 = imm_ujtype[19];
  assign _GEN_357 = csr__GEN_357_0;
  assign _GEN_160_0 = _T_306 | io_ctl_pipeline_kill;
  assign _GEN_279 = csr__GEN_279_0;
  assign _GEN_133_0 = ~io_ctl_full_stall;
  assign _GEN_399 = csr__GEN_399_0;
  assign _GEN_264 = csr__GEN_264_0;
  assign _GEN_300 = csr__GEN_300_0;
  assign _GEN_127_0 = _T_306 | io_ctl_pipeline_kill;
  assign _GEN_432 = csr__GEN_432_0;
  assign _GEN_381 = csr__GEN_381_0;
  assign _GEN_339_0 = csr__GEN_339_1;
  assign _GEN_261 = csr__GEN_261_0;
  assign _GEN_16_0 = io_ctl_exe_pc_sel == 2'h1;
  assign _GEN_360 = csr__GEN_360_0;
  assign _GEN_163_0 = reset;
  assign _GEN_246_0 = csr__GEN_246_1;
  assign _GEN_438 = csr__GEN_438_0;
  assign _GEN_282 = csr__GEN_282_0;
  assign _GEN_345_0 = csr__GEN_345_1;
  assign _GEN_121_0 = _T_145 & _T_147;
  assign _GEN_240_0 = csr__GEN_240_1;
  assign _GEN_148_0 = io_ctl_mem_exception;
  assign _GEN_154_0 = _T_306 | io_ctl_pipeline_kill;
  assign _GEN_444 = csr__GEN_444_0;
  assign _GEN_267_0 = csr__GEN_267_1;
  assign _GEN_459 = csr__GEN_459_0;
  assign _GEN_453 = csr__GEN_453_0;
  assign _GEN_366 = csr__GEN_366_0;
  assign _GEN_7_0 = csr__GEN_7_0;
  assign _GEN_142_0 = ~io_ctl_full_stall;
  assign _GEN_324_0 = csr__GEN_324_1;
  assign _GEN_333_0 = csr__GEN_333_1;
  assign _GEN_342 = csr__GEN_342_0;
  assign _GEN_405 = csr__GEN_405_0;
  assign _GEN_420_0 = csr__GEN_420_1;
  assign _GEN_306 = csr__GEN_306_0;
  assign _GEN_109_1 = _T_145 & _T_147;
  assign _GEN_103_0 = io_ctl_dec_kill;
  assign _GEN_3_0 = csr__GEN_3_0;
  assign _GEN_136_0 = ~io_ctl_full_stall;
  assign _GEN_426 = csr__GEN_426_0;
  assign _GEN_441 = csr__GEN_441_0;
  assign _GEN_94_1 = io_ctl_op1_sel == 2'h2;
  assign _GEN_348 = csr__GEN_348_0;
  assign _GEN_255 = csr__GEN_255_0;
  assign _GEN_115_0 = _T_145 & _T_147;
  assign _GEN_146_0 = csr__GEN_146_0;
  assign _GEN_363 = csr__GEN_363_0;
  assign _GEN_321_0 = csr__GEN_321_1;
  assign _GEN_327_0 = csr__GEN_327_1;
  assign _GEN_354 = csr__GEN_354_0;
  assign _GEN_234_0 = csr__GEN_234_1;
  assign _GEN_130_0 = _T_306 | io_ctl_pipeline_kill;
  assign _GEN_249_0 = csr__GEN_249_1;
  assign _GEN_243 = csr__GEN_243_0;
  assign _GEN_447 = csr__GEN_447_0;
  assign _GEN_330_0 = csr__GEN_330_1;
  assign _GEN_429 = csr__GEN_429_0;
  assign _GEN_293_0 = csr__GEN_293_1;
  assign _GEN_87_0 = exe_reg_ctrl_alu_fun == 4'h7;
  assign _GEN_414_0 = csr__GEN_414_1;
  assign _GEN_309 = csr__GEN_309_0;
  assign _GEN_299_0 = csr__GEN_299_1;
  assign _GEN_336 = csr__GEN_336_0;
  assign _GEN_408 = csr__GEN_408_0;
  assign _GEN_112_0 = _T_145 & _T_147;
  assign _GEN_150_0 = csr__GEN_150_0;
  assign _GEN_435 = csr__GEN_435_0;
  assign _GEN_97_1 = _T_266 & _T_224;
  assign _GEN_124_0 = _T_306 | io_ctl_pipeline_kill;
  assign _GEN_118_0 = _T_145 & _T_147;
  assign _GEN_392_0 = csr__GEN_392_1;
  assign _GEN_398_0 = csr__GEN_398_1;
  assign _GEN_423_0 = csr__GEN_423_1;
  assign _GEN_237 = csr__GEN_237_0;
  assign _GEN_315_0 = csr__GEN_315_1;
  assign _GEN_79_0 = exe_reg_ctrl_alu_fun == 4'ha;
  assign _GEN_1_2 = io_ctl_exe_pc_sel == 2'h2;
  assign _GEN_90_0 = exe_reg_ctrl_alu_fun == 4'h1;
  assign _GEN_162_0 = reset;
  assign _GEN_302_0 = csr__GEN_302_1;
  assign _GEN_106_1 = io_ctl_dec_kill;
  assign _GEN_71_1 = mem_reg_ctrl_wb_sel == 2'h3;
  assign _GEN_380_0 = csr__GEN_380_1;
  assign _GEN_174_0 = reset;
  assign _GEN_318_0 = csr__GEN_318_1;
  assign _GEN_287_0 = csr__GEN_287_1;
  assign _GEN_386_0 = csr__GEN_386_1;
  assign _GEN_281_0 = csr__GEN_281_1;
  assign _GEN_312_0 = csr__GEN_312_1;
  assign _GEN_417_0 = csr__GEN_417_1;
  assign _GEN_411_0 = csr__GEN_411_1;
  assign _GEN_55_1 = io_ctl_op2_sel == 3'h4;
  assign _GEN_100_1 = _T_265 & exe_reg_ctrl_rf_wen;
  assign _GEN_168_1 = io_ctl_pipeline_kill;
  assign _GEN_401_0 = csr__GEN_401_1;
  assign _GEN_44_1 = io_ctl_pipeline_kill;
  assign _GEN_74_1 = mem_reg_ctrl_wb_sel == 2'h0;
  assign _GEN_374_0 = csr__GEN_374_1;
  assign _GEN_368_0 = csr__GEN_368_1;
  assign _GEN_383_0 = csr__GEN_383_1;
  assign _GEN_263_0 = csr__GEN_263_1;
  assign _GEN_177_0 = ~io_ctl_full_stall;
  assign _GEN_171_0 = reset;
  assign _GEN_446 = csr__GEN_446_0;
  assign _GEN_290_0 = csr__GEN_290_1;
  assign _GEN_83_0 = exe_reg_ctrl_alu_fun == 4'h2;
  assign _GEN_135_1 = ~io_ctl_full_stall;
  assign _GEN_389_0 = csr__GEN_389_1;
  assign _GEN_93_0 = io_ctl_op1_sel == 2'h1;
  assign _GEN_254_0 = csr__GEN_254_1;
  assign _GEN_21_0 = _T_165 & _T_167;
  assign _GEN_461 = csr__GEN_461_0;
  assign _GEN_362_0 = csr__GEN_362_1;
  assign _GEN_156_0 = _T_306 | io_ctl_pipeline_kill;
  assign _GEN_150_1 = reset;
  assign _GEN_68_1 = io_ctl_op2_sel == 3'h1;
  assign _GEN_296_0 = csr__GEN_296_1;
  assign _GEN_395_0 = csr__GEN_395_1;
  assign _GEN_275_0 = csr__GEN_275_1;
  assign _GEN_269_0 = csr__GEN_269_1;
  assign _GEN_278_0 = csr__GEN_278_1;
  assign _GEN_138_0 = ~io_ctl_full_stall;
  assign _GEN_251_0 = csr__GEN_251_1;
  assign _GEN_455 = csr__GEN_455_0;
  assign _GEN_377_0 = csr__GEN_377_1;
  assign _GEN_153_1 = reset;
  assign _GEN_272_0 = csr__GEN_272_1;
  assign _GEN_47_1 = imm_sbtype[11];
  assign _GEN_335_0 = csr__GEN_335_1;
  assign _GEN_41_1 = _T_145 & _T_147;
  assign _GEN_434 = csr__GEN_434_0;
  assign _GEN_257_0 = csr__GEN_257_1;
  assign _GEN_443 = csr__GEN_443_0;
  assign _GEN_356_0 = csr__GEN_356_1;
  assign _GEN_350_0 = csr__GEN_350_1;
  assign _GEN_132_1 = ~io_ctl_full_stall;
  assign _GEN_144_0 = io_ctl_pipeline_kill;
  assign _GEN_159_0 = _T_306 | io_ctl_pipeline_kill;
  assign _GEN_428 = csr__GEN_428_0;
  assign _GEN_449 = csr__GEN_449_0;
  assign _GEN_117_1 = _T_145 & _T_147;
  assign _GEN_236_0 = csr__GEN_236_1;
  assign _GEN_371_0 = csr__GEN_371_1;
  assign _GEN_165_0 = reset;
  assign _GEN_284_0 = csr__GEN_284_1;
  assign _GEN_147_1 = io_ctl_pipeline_kill;
  assign _GEN_416_0 = csr__GEN_416_1;
  assign _GEN_260_0 = csr__GEN_260_1;
  assign _GEN_105_1 = io_ctl_dec_kill;
  assign _GEN_338_0 = csr__GEN_338_1;
  assign _GEN_141_1 = ~io_ctl_full_stall;
  assign _GEN_99_1 = _T_272 & mem_reg_ctrl_rf_wen;
  assign _GEN_344_0 = csr__GEN_344_1;
  assign _GEN_239_0 = csr__GEN_239_1;
  assign _GEN_353_0 = csr__GEN_353_1;
  assign _GEN_266_0 = csr__GEN_266_1;
  assign _GEN_452 = csr__GEN_452_0;
  assign _GEN_120_1 = _T_145 & _T_147;
  assign _GEN_365_0 = csr__GEN_365_1;
  assign _GEN_6_0 = csr__GEN_6_0;
  assign _GEN_410_0 = csr__GEN_410_1;
  assign _GEN_152_1 = csr__GEN_152_1;
  assign _GEN_437 = csr__GEN_437_0;
  assign _GEN_332_0 = csr__GEN_332_1;
  assign _GEN_126_1 = _T_306 | io_ctl_pipeline_kill;
  assign _GEN_245_0 = csr__GEN_245_1;
  assign _GEN_359_0 = csr__GEN_359_1;
  assign _GEN_431 = csr__GEN_431_0;
  assign _GEN_458 = csr__GEN_458_0;
  assign _GEN_317_0 = csr__GEN_317_1;
  assign _GEN_326_0 = csr__GEN_326_1;
  assign _GEN_341_0 = csr__GEN_341_1;
  assign _GEN_1_3 = regfile__GEN_1_3;
  assign _GEN_394_0 = csr__GEN_394_1;
  assign _GEN_248_0 = csr__GEN_248_1;
  assign _GEN_347_0 = csr__GEN_347_1;
  assign _GEN_92_1 = _T_245 & exe_reg_ctrl_rf_wen;
  assign _GEN_102_1 = io_ctl_dec_kill;
  assign _GEN_425_0 = csr__GEN_425_1;
  assign _GEN_305_0 = csr__GEN_305_1;
  assign _GEN_419_0 = csr__GEN_419_1;
  assign _GEN_320_0 = csr__GEN_320_1;
  assign _GEN_108_1 = io_ctl_dec_kill;
  assign _GEN_114_1 = _T_145 & _T_147;
  assign _GEN_123_1 = _T_306 | io_ctl_pipeline_kill;
  assign _GEN_413_0 = csr__GEN_413_1;
  assign _GEN_440 = csr__GEN_440_0;
  assign _GEN_295_0 = csr__GEN_295_1;
  assign _GEN_129_1 = _T_306 | io_ctl_pipeline_kill;
  assign _GEN_404_0 = csr__GEN_404_1;
  assign _GEN_403_0 = csr__GEN_403_1;
  assign _GEN_242_0 = csr__GEN_242_1;
  assign _GEN_15_1 = csr__GEN_15_1;
  assign _GEN_96_1 = _T_273 & _T_224;
  assign _GEN_86_1 = exe_reg_ctrl_alu_fun == 4'h8;
  assign _GEN_164_1 = reset;
  assign _GEN_308_0 = csr__GEN_308_1;
  assign _GEN_149_1 = csr__GEN_149_1;
  assign _GEN_329_0 = csr__GEN_329_1;
  assign _GEN_292_0 = csr__GEN_292_1;
  assign _GEN_298_0 = csr__GEN_298_1;
  assign _GEN_391_0 = csr__GEN_391_1;
  assign _GEN_314_0 = csr__GEN_314_1;
  assign _GEN_323_0 = csr__GEN_323_1;
  assign _GEN_376_0 = csr__GEN_376_1;
  assign _GEN_422_0 = csr__GEN_422_1;
  assign _GEN_277_0 = csr__GEN_277_1;
  assign _GEN_46_1 = imm_stype[11];
  assign _GEN_111_1 = _T_145 & _T_147;
  assign _GEN_78_1 = exe_reg_ctrl_alu_fun == 4'hb;
  assign _GEN_407_0 = csr__GEN_407_1;
  assign _GEN_179_1 = reset;
  assign _GEN_397_0 = csr__GEN_397_1;
  assign _GEN_173_1 = reset;
  assign _GEN_70_1 = _T_255 & wb_reg_ctrl_rf_wen;
  assign _GEN_379_0 = csr__GEN_379_1;
  assign _GEN_82_1 = exe_reg_ctrl_alu_fun == 4'h4;
  assign _GEN_373_0 = csr__GEN_373_1;
  assign _GEN_54_1 = io_ctl_op2_sel == 3'h5;
  assign _GEN_364_0 = csr__GEN_364_1;
  assign _GEN_259_0 = csr__GEN_259_1;
  assign _GEN_167_1 = io_ctl_pipeline_kill;
  assign _GEN_43_1 = io_ctl_pipeline_kill;
  assign _GEN_161_1 = reset;
  assign _GEN_265_0 = csr__GEN_265_1;
  assign _GEN_301_0 = csr__GEN_301_1;
  assign _GEN_146_2 = io_ctl_pipeline_kill;
  assign _GEN_286_0 = csr__GEN_286_1;
  assign _GEN_400_0 = csr__GEN_400_1;
  assign _GEN_89_0 = exe_reg_ctrl_alu_fun == 4'h5;
  assign _GEN_358_0 = csr__GEN_358_1;
  assign _GEN_385_0 = csr__GEN_385_1;
  assign _GEN_457 = csr__GEN_457_0;
  assign _GEN_311_0 = csr__GEN_311_1;
  assign _GEN_280_0 = csr__GEN_280_1;
  assign _GEN_143_1 = io_ctl_pipeline_kill;
  assign _GEN_367_0 = csr__GEN_367_1;
  assign _GEN_247_0 = csr__GEN_247_1;
  assign _GEN_274_0 = csr__GEN_274_1;
  assign _GEN_460 = csr__GEN_460_0;
  assign _GEN_283_0 = csr__GEN_283_1;
  assign _GEN_388_0 = csr__GEN_388_1;
  assign _GEN_382_0 = csr__GEN_382_1;
  assign _GEN_268_0 = csr__GEN_268_1;
  assign _GEN_176_1 = reset;
  assign _GEN_346_0 = csr__GEN_346_1;
  assign _GEN_64_1 = io_ctl_op2_sel == 3'h2;
  assign _GEN_340_0 = csr__GEN_340_1;
  assign _GEN_134_1 = ~io_ctl_full_stall;
  assign _GEN_149_2 = reset;
  assign _GEN_439 = csr__GEN_439_0;
  assign _GEN_262_0 = csr__GEN_262_1;
  assign _GEN_17_1 = io_ctl_exe_pc_sel == 2'h0;
  assign _GEN_361_0 = csr__GEN_361_1;
  assign _GEN_155_1 = _T_306 | io_ctl_pipeline_kill;
  assign _GEN_170_1 = io_ctl_pipeline_kill;
  assign _GEN_73_1 = mem_reg_ctrl_wb_sel == 2'h2;
  assign _GEN_128_1 = _T_306 | io_ctl_pipeline_kill;
  assign _GEN_241_0 = csr__GEN_241_1;
  assign _GEN_445 = csr__GEN_445_0;
  assign _GEN_289_0 = csr__GEN_289_1;
  assign _GEN_131_1 = exe_reg_ctrl_wb_sel == 2'h2;
  assign _GEN_152_2 = reset;
  assign _GEN_421_0 = csr__GEN_421_1;
  assign _GEN_427 = csr__GEN_427_0;
  assign _GEN_454 = csr__GEN_454_0;
  assign _GEN_256_0 = csr__GEN_256_1;
  assign _GEN_110_1 = _T_145 & _T_147;
  assign _GEN_40_1 = io_ctl_if_kill;
  assign _GEN_5_2 = csr__GEN_5_2;
  assign _GEN_158_1 = reset;
  assign _GEN_271_0 = csr__GEN_271_1;
  assign _GEN_322_0 = csr__GEN_322_1;
  assign _GEN_334_0 = csr__GEN_334_1;
  assign _GEN_116_1 = _T_145 & _T_147;
  assign _GEN_235_0 = csr__GEN_235_1;
  assign _GEN_349_0 = csr__GEN_349_1;
  assign _GEN_147_2 = csr__GEN_147_2;
  assign _GEN_448 = csr__GEN_448_0;
  assign _GEN_442 = csr__GEN_442_0;
  assign _GEN_343_0 = csr__GEN_343_1;
  assign _GEN_355_0 = csr__GEN_355_1;
  assign _GEN_137_1 = ~io_ctl_full_stall;
  assign _GEN_370_0 = csr__GEN_370_1;
  assign _GEN_250_0 = csr__GEN_250_1;
  assign _GEN_463 = csr__GEN_463_0;
  assign _GEN_328_0 = csr__GEN_328_1;
  assign regfile_clock = clock;
  assign regfile_io_rs1_addr = dec_reg_inst[19:15]; // @[dpath.scala 158:24]
  assign regfile_io_rs2_addr = dec_reg_inst[24:20]; // @[dpath.scala 159:24]
  assign regfile_io_waddr = wb_reg_wbaddr; // @[dpath.scala 162:21]
  assign regfile_io_wdata = wb_reg_wbdata; // @[dpath.scala 163:21]
  assign regfile_io_wen = wb_reg_ctrl_rf_wen; // @[dpath.scala 164:21]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_rw_cmd = mem_reg_ctrl_csr_cmd; // @[dpath.scala 360:20]
  assign csr_io_rw_wdata = mem_reg_alu_out; // @[dpath.scala 359:20]
  assign csr_io_decode_csr = mem_reg_inst[31:20]; // @[dpath.scala 358:23]
  assign csr_io_exception = io_ctl_mem_exception; // @[dpath.scala 363:21]
  assign csr_io_retire = _T_147 & _T_145; // @[dpath.scala 362:21]
  assign csr_io_pc = mem_reg_pc; // @[dpath.scala 364:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  if_reg_pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  dec_reg_inst = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  dec_reg_pc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  exe_reg_inst = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  exe_reg_pc = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  exe_reg_wbaddr = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  exe_alu_op1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  brjmp_offset = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  exe_reg_rs2_data = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  exe_reg_ctrl_br_type = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  exe_reg_ctrl_alu_fun = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  exe_reg_ctrl_wb_sel = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  exe_reg_ctrl_rf_wen = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  exe_reg_ctrl_mem_val = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  exe_reg_ctrl_mem_fcn = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  exe_reg_ctrl_mem_typ = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  exe_reg_ctrl_csr_cmd = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  mem_reg_pc = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  mem_reg_inst = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  mem_reg_alu_out = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  mem_reg_wbaddr = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  mem_reg_rs2_data = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  mem_reg_ctrl_rf_wen = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  mem_reg_ctrl_mem_val = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  mem_reg_ctrl_mem_fcn = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  mem_reg_ctrl_mem_typ = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  mem_reg_ctrl_wb_sel = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  mem_reg_ctrl_csr_cmd = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  wb_reg_wbaddr = _RAND_28[4:0];
  _RAND_29 = {1{`RANDOM}};
  wb_reg_wbdata = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  wb_reg_ctrl_rf_wen = _RAND_30[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      if_reg_pc <= 32'h0;
    end else if (reset) begin
      if_reg_pc <= 32'h80000000;
    end else if (_T_149) begin
      if (!(_T_168)) begin
        if (_T_158) begin
          if_reg_pc <= if_pc_plus4;
        end else if (_T_153) begin
          if_reg_pc <= exe_brjmp_target;
        end else if (_T_154) begin
          if_reg_pc <= exe_adder_out;
        end else begin
          if_reg_pc <= exception_target;
        end
      end
    end
    if (metaReset) begin
      dec_reg_inst <= 32'h0;
    end else if (reset) begin
      dec_reg_inst <= 32'h4033;
    end else if (io_ctl_pipeline_kill) begin
      dec_reg_inst <= 32'h4033;
    end else if (_T_148) begin
      if (io_ctl_if_kill) begin
        dec_reg_inst <= 32'h4033;
      end else begin
        dec_reg_inst <= io_imem_resp_bits_data;
      end
    end
    if (metaReset) begin
      dec_reg_pc <= 32'h0;
    end else if (reset) begin
      dec_reg_pc <= 32'h0;
    end else if (!(io_ctl_pipeline_kill)) begin
      if (_T_148) begin
        dec_reg_pc <= if_reg_pc;
      end
    end
    if (metaReset) begin
      exe_reg_inst <= 32'h0;
    end else if (reset) begin
      exe_reg_inst <= 32'h4033;
    end else if (_T_307) begin
      exe_reg_inst <= 32'h4033;
    end else if (_T_148) begin
      if (io_ctl_dec_kill) begin
        exe_reg_inst <= 32'h4033;
      end else begin
        exe_reg_inst <= dec_reg_inst;
      end
    end
    if (metaReset) begin
      exe_reg_pc <= 32'h0;
    end else if (reset) begin
      exe_reg_pc <= 32'h0;
    end else if (!(_T_307)) begin
      if (_T_148) begin
        exe_reg_pc <= dec_reg_pc;
      end
    end
    if (metaReset) begin
      exe_reg_wbaddr <= 5'h0;
    end else if (_T_307) begin
      exe_reg_wbaddr <= 5'h0;
    end else if (_T_148) begin
      if (io_ctl_dec_kill) begin
        exe_reg_wbaddr <= 5'h0;
      end else begin
        exe_reg_wbaddr <= dec_wbaddr;
      end
    end
    if (metaReset) begin
      exe_alu_op1 <= 32'h0;
    end else if (!(_T_307)) begin
      if (_T_148) begin
        if (_T_240) begin
          exe_alu_op1 <= imm_z;
        end else if (_T_241) begin
          exe_alu_op1 <= dec_reg_pc;
        end else if (_T_246) begin
          if (_T_321) begin
            exe_alu_op1 <= exe_adder_out;
          end else if (_T_322) begin
            exe_alu_op1 <= _T_325;
          end else if (_T_326) begin
            exe_alu_op1 <= _T_327;
          end else if (_T_328) begin
            exe_alu_op1 <= _T_329;
          end else if (_T_330) begin
            exe_alu_op1 <= _T_331;
          end else if (_T_332) begin
            exe_alu_op1 <= {{31'd0}, _T_335};
          end else if (_T_336) begin
            exe_alu_op1 <= {{31'd0}, _T_337};
          end else if (_T_338) begin
            exe_alu_op1 <= _T_339[31:0];
          end else if (_T_341) begin
            exe_alu_op1 <= _T_344;
          end else if (_T_345) begin
            exe_alu_op1 <= _T_346;
          end else if (!(_T_347)) begin
            if (_T_348) begin
              exe_alu_op1 <= brjmp_offset;
            end else begin
              exe_alu_op1 <= exe_reg_inst;
            end
          end
        end else if (_T_251) begin
          if (_T_439) begin
            exe_alu_op1 <= mem_reg_alu_out;
          end else if (_T_440) begin
            exe_alu_op1 <= mem_reg_alu_out;
          end else if (_T_441) begin
            exe_alu_op1 <= io_dmem_resp_bits_data;
          end else if (_T_442) begin
            exe_alu_op1 <= csr_io_rw_rdata;
          end else begin
            exe_alu_op1 <= mem_reg_alu_out;
          end
        end else if (_T_256) begin
          exe_alu_op1 <= wb_reg_wbdata;
        end else begin
          exe_alu_op1 <= regfile_io_rs1_data;
        end
      end
    end
    if (metaReset) begin
      brjmp_offset <= 32'h0;
    end else if (!(_T_307)) begin
      if (_T_148) begin
        if (_T_268) begin
          if (_T_321) begin
            brjmp_offset <= exe_adder_out;
          end else if (_T_322) begin
            brjmp_offset <= _T_325;
          end else if (_T_326) begin
            brjmp_offset <= _T_327;
          end else if (_T_328) begin
            brjmp_offset <= _T_329;
          end else if (_T_330) begin
            brjmp_offset <= _T_331;
          end else if (_T_332) begin
            brjmp_offset <= {{31'd0}, _T_335};
          end else if (_T_336) begin
            brjmp_offset <= {{31'd0}, _T_337};
          end else if (_T_338) begin
            brjmp_offset <= _T_339[31:0];
          end else if (_T_341) begin
            brjmp_offset <= _T_344;
          end else if (_T_345) begin
            brjmp_offset <= _T_346;
          end else if (_T_347) begin
            brjmp_offset <= exe_alu_op1;
          end else if (!(_T_348)) begin
            brjmp_offset <= exe_reg_inst;
          end
        end else if (_T_275) begin
          if (_T_439) begin
            brjmp_offset <= mem_reg_alu_out;
          end else if (_T_440) begin
            brjmp_offset <= mem_reg_alu_out;
          end else if (_T_441) begin
            brjmp_offset <= io_dmem_resp_bits_data;
          end else if (_T_442) begin
            brjmp_offset <= csr_io_rw_rdata;
          end else begin
            brjmp_offset <= mem_reg_alu_out;
          end
        end else if (_T_282) begin
          brjmp_offset <= wb_reg_wbdata;
        end else if (_T_224) begin
          brjmp_offset <= regfile_io_rs2_data;
        end else if (_T_225) begin
          brjmp_offset <= imm_itype_sext;
        end else if (_T_226) begin
          brjmp_offset <= imm_stype_sext;
        end else if (_T_227) begin
          brjmp_offset <= imm_sbtype_sext;
        end else if (_T_228) begin
          brjmp_offset <= imm_utype_sext;
        end else if (_T_229) begin
          brjmp_offset <= imm_ujtype_sext;
        end else begin
          brjmp_offset <= 32'h0;
        end
      end
    end
    if (metaReset) begin
      exe_reg_rs2_data <= 32'h0;
    end else if (!(_T_307)) begin
      if (_T_148) begin
        if (_T_266) begin
          if (_T_321) begin
            exe_reg_rs2_data <= exe_adder_out;
          end else if (_T_322) begin
            exe_reg_rs2_data <= _T_325;
          end else if (_T_326) begin
            exe_reg_rs2_data <= _T_327;
          end else if (_T_328) begin
            exe_reg_rs2_data <= _T_329;
          end else if (_T_330) begin
            exe_reg_rs2_data <= _T_331;
          end else if (_T_332) begin
            exe_reg_rs2_data <= {{31'd0}, _T_335};
          end else if (_T_336) begin
            exe_reg_rs2_data <= {{31'd0}, _T_337};
          end else if (_T_338) begin
            exe_reg_rs2_data <= _T_339[31:0];
          end else if (_T_341) begin
            exe_reg_rs2_data <= _T_344;
          end else if (_T_345) begin
            exe_reg_rs2_data <= _T_346;
          end else if (_T_347) begin
            exe_reg_rs2_data <= exe_alu_op1;
          end else if (_T_348) begin
            exe_reg_rs2_data <= brjmp_offset;
          end else begin
            exe_reg_rs2_data <= exe_reg_inst;
          end
        end else if (_T_273) begin
          if (_T_439) begin
            exe_reg_rs2_data <= mem_reg_alu_out;
          end else if (_T_440) begin
            exe_reg_rs2_data <= mem_reg_alu_out;
          end else if (_T_441) begin
            exe_reg_rs2_data <= io_dmem_resp_bits_data;
          end else if (_T_442) begin
            exe_reg_rs2_data <= csr_io_rw_rdata;
          end else begin
            exe_reg_rs2_data <= mem_reg_alu_out;
          end
        end else if (_T_280) begin
          exe_reg_rs2_data <= wb_reg_wbdata;
        end else begin
          exe_reg_rs2_data <= regfile_io_rs2_data;
        end
      end
    end
    if (metaReset) begin
      exe_reg_ctrl_br_type <= 4'h0;
    end else if (reset) begin
      exe_reg_ctrl_br_type <= 4'h0;
    end else if (_T_307) begin
      exe_reg_ctrl_br_type <= 4'h0;
    end else if (_T_148) begin
      if (io_ctl_dec_kill) begin
        exe_reg_ctrl_br_type <= 4'h0;
      end else begin
        exe_reg_ctrl_br_type <= io_ctl_br_type;
      end
    end
    if (metaReset) begin
      exe_reg_ctrl_alu_fun <= 4'h0;
    end else if (!(_T_307)) begin
      if (_T_148) begin
        exe_reg_ctrl_alu_fun <= io_ctl_alu_fun;
      end
    end
    if (metaReset) begin
      exe_reg_ctrl_wb_sel <= 2'h0;
    end else if (!(_T_307)) begin
      if (_T_148) begin
        exe_reg_ctrl_wb_sel <= io_ctl_wb_sel;
      end
    end
    if (metaReset) begin
      exe_reg_ctrl_rf_wen <= 1'h0;
    end else if (reset) begin
      exe_reg_ctrl_rf_wen <= 1'h0;
    end else if (_T_307) begin
      exe_reg_ctrl_rf_wen <= 1'h0;
    end else if (_T_148) begin
      if (io_ctl_dec_kill) begin
        exe_reg_ctrl_rf_wen <= 1'h0;
      end else begin
        exe_reg_ctrl_rf_wen <= io_ctl_rf_wen;
      end
    end
    if (metaReset) begin
      exe_reg_ctrl_mem_val <= 1'h0;
    end else if (reset) begin
      exe_reg_ctrl_mem_val <= 1'h0;
    end else if (_T_307) begin
      exe_reg_ctrl_mem_val <= 1'h0;
    end else if (_T_148) begin
      if (io_ctl_dec_kill) begin
        exe_reg_ctrl_mem_val <= 1'h0;
      end else begin
        exe_reg_ctrl_mem_val <= io_ctl_mem_val;
      end
    end
    if (metaReset) begin
      exe_reg_ctrl_mem_fcn <= 1'h0;
    end else if (reset) begin
      exe_reg_ctrl_mem_fcn <= 1'h0;
    end else begin
      exe_reg_ctrl_mem_fcn <= _GEN_36[0];
    end
    if (metaReset) begin
      exe_reg_ctrl_mem_typ <= 3'h0;
    end else if (reset) begin
      exe_reg_ctrl_mem_typ <= 3'h0;
    end else if (!(_T_307)) begin
      if (_T_148) begin
        if (!(io_ctl_dec_kill)) begin
          exe_reg_ctrl_mem_typ <= io_ctl_mem_typ;
        end
      end
    end
    if (metaReset) begin
      exe_reg_ctrl_csr_cmd <= 3'h0;
    end else if (reset) begin
      exe_reg_ctrl_csr_cmd <= 3'h0;
    end else if (_T_307) begin
      exe_reg_ctrl_csr_cmd <= 3'h0;
    end else if (_T_148) begin
      if (io_ctl_dec_kill) begin
        exe_reg_ctrl_csr_cmd <= 3'h0;
      end else begin
        exe_reg_ctrl_csr_cmd <= io_ctl_csr_cmd;
      end
    end
    if (metaReset) begin
      mem_reg_pc <= 32'h0;
    end else if (io_ctl_pipeline_kill) begin
      mem_reg_pc <= 32'h4033;
    end else if (_T_147) begin
      mem_reg_pc <= exe_reg_pc;
    end
    if (metaReset) begin
      mem_reg_inst <= 32'h0;
    end else if (!(io_ctl_pipeline_kill)) begin
      if (_T_147) begin
        mem_reg_inst <= exe_reg_inst;
      end
    end
    if (metaReset) begin
      mem_reg_alu_out <= 32'h0;
    end else if (!(io_ctl_pipeline_kill)) begin
      if (_T_147) begin
        if (_T_371) begin
          mem_reg_alu_out <= exe_pc_plus4;
        end else if (_T_321) begin
          mem_reg_alu_out <= exe_adder_out;
        end else if (_T_322) begin
          mem_reg_alu_out <= _T_325;
        end else if (_T_326) begin
          mem_reg_alu_out <= _T_327;
        end else if (_T_328) begin
          mem_reg_alu_out <= _T_329;
        end else if (_T_330) begin
          mem_reg_alu_out <= _T_331;
        end else if (_T_332) begin
          mem_reg_alu_out <= {{31'd0}, _T_335};
        end else if (_T_336) begin
          mem_reg_alu_out <= {{31'd0}, _T_337};
        end else if (_T_338) begin
          mem_reg_alu_out <= _T_339[31:0];
        end else if (_T_341) begin
          mem_reg_alu_out <= _T_344;
        end else if (_T_345) begin
          mem_reg_alu_out <= _T_346;
        end else if (_T_347) begin
          mem_reg_alu_out <= exe_alu_op1;
        end else if (_T_348) begin
          mem_reg_alu_out <= brjmp_offset;
        end else begin
          mem_reg_alu_out <= exe_reg_inst;
        end
      end
    end
    if (metaReset) begin
      mem_reg_wbaddr <= 5'h0;
    end else if (!(io_ctl_pipeline_kill)) begin
      if (_T_147) begin
        mem_reg_wbaddr <= exe_reg_wbaddr;
      end
    end
    if (metaReset) begin
      mem_reg_rs2_data <= 32'h0;
    end else if (!(io_ctl_pipeline_kill)) begin
      if (_T_147) begin
        mem_reg_rs2_data <= exe_reg_rs2_data;
      end
    end
    if (metaReset) begin
      mem_reg_ctrl_rf_wen <= 1'h0;
    end else if (reset) begin
      mem_reg_ctrl_rf_wen <= 1'h0;
    end else if (io_ctl_pipeline_kill) begin
      mem_reg_ctrl_rf_wen <= 1'h0;
    end else if (_T_147) begin
      mem_reg_ctrl_rf_wen <= exe_reg_ctrl_rf_wen;
    end
    if (metaReset) begin
      mem_reg_ctrl_mem_val <= 1'h0;
    end else if (reset) begin
      mem_reg_ctrl_mem_val <= 1'h0;
    end else if (io_ctl_pipeline_kill) begin
      mem_reg_ctrl_mem_val <= 1'h0;
    end else if (_T_147) begin
      mem_reg_ctrl_mem_val <= exe_reg_ctrl_mem_val;
    end
    if (metaReset) begin
      mem_reg_ctrl_mem_fcn <= 1'h0;
    end else if (reset) begin
      mem_reg_ctrl_mem_fcn <= 1'h0;
    end else if (!(io_ctl_pipeline_kill)) begin
      if (_T_147) begin
        mem_reg_ctrl_mem_fcn <= exe_reg_ctrl_mem_fcn;
      end
    end
    if (metaReset) begin
      mem_reg_ctrl_mem_typ <= 3'h0;
    end else if (reset) begin
      mem_reg_ctrl_mem_typ <= 3'h0;
    end else if (!(io_ctl_pipeline_kill)) begin
      if (_T_147) begin
        mem_reg_ctrl_mem_typ <= exe_reg_ctrl_mem_typ;
      end
    end
    if (metaReset) begin
      mem_reg_ctrl_wb_sel <= 2'h0;
    end else if (!(io_ctl_pipeline_kill)) begin
      if (_T_147) begin
        mem_reg_ctrl_wb_sel <= exe_reg_ctrl_wb_sel;
      end
    end
    if (metaReset) begin
      mem_reg_ctrl_csr_cmd <= 3'h0;
    end else if (reset) begin
      mem_reg_ctrl_csr_cmd <= 3'h0;
    end else if (io_ctl_pipeline_kill) begin
      mem_reg_ctrl_csr_cmd <= 3'h0;
    end else if (_T_147) begin
      mem_reg_ctrl_csr_cmd <= exe_reg_ctrl_csr_cmd;
    end
    if (metaReset) begin
      wb_reg_wbaddr <= 5'h0;
    end else if (_T_147) begin
      wb_reg_wbaddr <= mem_reg_wbaddr;
    end
    if (metaReset) begin
      wb_reg_wbdata <= 32'h0;
    end else if (_T_147) begin
      if (_T_439) begin
        wb_reg_wbdata <= mem_reg_alu_out;
      end else if (_T_440) begin
        wb_reg_wbdata <= mem_reg_alu_out;
      end else if (_T_441) begin
        wb_reg_wbdata <= io_dmem_resp_bits_data;
      end else if (_T_442) begin
        wb_reg_wbdata <= csr_io_rw_rdata;
      end else begin
        wb_reg_wbdata <= mem_reg_alu_out;
      end
    end
    if (metaReset) begin
      wb_reg_ctrl_rf_wen <= 1'h0;
    end else if (reset) begin
      wb_reg_ctrl_rf_wen <= 1'h0;
    end else begin
      wb_reg_ctrl_rf_wen <= _GEN_81;
    end
  end
endmodule
module Core(
  input         metaReset,
  input         clock,
  input         reset,
  output [31:0] io_imem_req_bits_addr,
  input         io_imem_resp_valid,
  input  [31:0] io_imem_resp_bits_data,
  output        io_dmem_req_valid,
  output [31:0] io_dmem_req_bits_addr,
  output [31:0] io_dmem_req_bits_data,
  output        io_dmem_req_bits_fcn,
  output [2:0]  io_dmem_req_bits_typ,
  input         io_dmem_resp_valid,
  input  [31:0] io_dmem_resp_bits_data,
  output        _GEN_451,
  output        _GEN_331,
  output        _GEN_337,
  output        _GEN_113,
  output        _GEN_111,
  output        _GEN_415,
  output        _GEN_436,
  output        _GEN_140,
  output        _GEN_71,
  output        _GEN_324,
  output        _GEN_219,
  output        _GEN_168,
  output        _GEN_98,
  output        _GEN_1,
  output        _GEN_352,
  output        _GEN_423,
  output        _GEN_44,
  output        _GEN_125,
  output        _GEN_267,
  output        _GEN_126,
  output        _GEN_430,
  output        _GEN_153,
  output        _GEN_225,
  output        _GEN_119,
  output        _GEN_88,
  output        _GEN_59,
  output        _GEN_252,
  output        _GEN_151,
  output        _GEN_147,
  output        _GEN_310,
  output        _GEN_351,
  output        _GEN_210,
  output        _GEN_246,
  output        _GEN_104,
  output        _GEN_409,
  output        _GEN_65,
  output        _GEN_253,
  output        _GEN_132,
  output        _GEN_318,
  output        _GEN_316,
  output        _GEN_92,
  output        _GEN_345,
  output        _GEN_231,
  output        _GEN_417,
  output        _GEN_244,
  output        _GEN_50,
  output        _GEN_238,
  output        _GEN_330,
  output        _GEN_86,
  output        _GEN_339,
  output        _GEN_101,
  output        _GEN_325,
  output        _GEN_240,
  output        _GEN_234,
  output        _GEN_120,
  output        _GEN_169,
  output        _GEN_129,
  output        _GEN_433,
  output        _GEN_333,
  output        _GEN_302,
  output        _GEN_313,
  output        _GEN_228,
  output        _GEN_197,
  output        _GEN_91,
  output        _GEN_411,
  output        _GEN_11,
  output        _GEN_401,
  output        _GEN_47,
  output        _GEN_296,
  output        _GEN_304,
  output        _GEN_294,
  output        _GEN_74,
  output        _GEN_213,
  output        _GEN_303,
  output        _GEN_107,
  output        _GEN_32,
  output        _GEN_0,
  output        _GEN_402,
  output        _GEN_412,
  output        _GEN_68,
  output        _GEN_135,
  output        _GEN_424,
  output        _GEN_175,
  output        _GEN_319,
  output        _GEN_288,
  output        _GEN_56,
  output        _GEN_26,
  output        _GEN_418,
  output        _GEN_122,
  output        _GEN_387,
  output        _GEN_53,
  output        _GEN_141,
  output        _GEN_327,
  output        _GEN_72,
  output        _GEN_395,
  output        _GEN_249,
  output        _GEN_114,
  output        _GEN_312,
  output        _GEN_203,
  output        _GEN_75,
  output        _GEN_85,
  output        _GEN_20,
  output        _GEN_178,
  output        _GEN_15,
  output        _GEN_157,
  output        _GEN_462,
  output        _GEN_69,
  output        _GEN_216,
  output        _GEN_206,
  output        _GEN_375,
  output        _GEN_151_0,
  output        _GEN_420,
  output        _GEN_123,
  output        _GEN_315,
  output        _GEN_284,
  output        _GEN_179,
  output        _GEN_33,
  output        _GEN_222,
  output        _GEN_377,
  output        _GEN_191,
  output        _GEN_290,
  output        _GEN_404,
  output        _GEN_390,
  output        _GEN_56_0,
  output        _GEN_305,
  output        _GEN_299,
  output        _GEN_185,
  output        _GEN_307,
  output        _GEN_297,
  output        _GEN_398,
  output        _GEN_406,
  output        _GEN_41,
  output        _GEN_321,
  output        _GEN_270,
  output        _GEN_95,
  output        _GEN_45,
  output        _GEN_414,
  output        _GEN_383,
  output        _GEN_369,
  output        _GEN_35,
  output        _GEN_29,
  output        _GEN_278,
  output        _GEN_117,
  output        _GEN_396,
  output        _GEN_172,
  output        _GEN_276,
  output        _GEN_291,
  output        _GEN_365,
  output        _GEN_359,
  output        _GEN_258,
  output        _GEN_372,
  output        _GEN_38,
  output        _GEN_252_0,
  output        _GEN_167,
  output        _GEN_166,
  output        _GEN_285,
  output        _GEN_42,
  output        _GEN_350,
  output        _GEN_106,
  output        _GEN_384,
  output        _GEN_18,
  output        _GEN_378,
  output        _GEN_393,
  output        _GEN_273,
  output        _GEN_293,
  output        _GEN_456,
  output        _GEN_371,
  output        _GEN_80,
  output        _GEN_351_0,
  output        _GEN_251,
  output        _GEN_209,
  output        _GEN_139,
  output        _GEN_145,
  output        _GEN_450,
  output        _GEN_308,
  output        _GEN_173,
  output        _GEN_53_0,
  output        _GEN_357,
  output        _GEN_200,
  output        _GEN_386,
  output        _GEN_272,
  output        _GEN_160,
  output        _GEN_91_0,
  output        _GEN_279,
  output        _GEN_194,
  output        _GEN_188,
  output        _GEN_133,
  output        _GEN_392,
  output        _GEN_23,
  output        _GEN_407,
  output        _GEN_287,
  output        _GEN_266,
  output        _GEN_399,
  output        _GEN_264,
  output        _GEN_300,
  output        _GEN_374,
  output        _GEN_233,
  output        _GEN_127,
  output        _GEN_269,
  output        _GEN_432,
  output        _GEN_381,
  output        _GEN_260,
  output        _GEN_161,
  output        _GEN_155,
  output        _GEN_339_0,
  output        _GEN_368,
  output        _GEN_254,
  output        _GEN_281,
  output        _GEN_73,
  output        _GEN_261,
  output        _GEN_353,
  output        _GEN_332,
  output        _GEN_88_0,
  output        _GEN_176,
  output        _GEN_16,
  output        _GEN_380,
  output        _GEN_360,
  output        _GEN_389,
  output        _GEN_163,
  output        _GEN_246_0,
  output        _GEN_438,
  output        _GEN_94,
  output        _GEN_282,
  output        _GEN_347,
  output        _GEN_109,
  output        _GEN_182,
  output        _GEN_345_0,
  output        _GEN_121,
  output        _GEN_240_0,
  output        _GEN_9,
  output        _GEN_148,
  output        _GEN_154,
  output        _GEN_444,
  output        _GEN_149,
  output        _GEN_267_0,
  output        _GEN_459,
  output        _GEN_453,
  output        _GEN_248,
  output        _GEN_366,
  output        _GEN_7,
  output        _GEN_142,
  output        _GEN_275,
  output        _GEN_140_0,
  output        _GEN_324_0,
  output        _GEN_100,
  output        _GEN_333_0,
  output        _GEN_362,
  output        _GEN_413,
  output        _GEN_342,
  output        _GEN_405,
  output        _GEN_420_0,
  output        _GEN_306,
  output        _GEN_76,
  output        _GEN_164,
  output        _GEN_109_0,
  output        _GEN_103,
  output        _GEN_3,
  output        _GEN_242,
  output        _GEN_136,
  output        _GEN_426,
  output        _GEN_137,
  output        _GEN_441,
  output        _GEN_341,
  output        _GEN_94_0,
  output        _GEN_348,
  output        _GEN_263,
  output        _GEN_257,
  output        _GEN_122_0,
  output        _GEN_143,
  output        _GEN_255,
  output        _GEN_82,
  output        _GEN_170,
  output        _GEN_356,
  output        _GEN_221,
  output        _GEN_215,
  output        _GEN_115,
  output        _GEN_146,
  output        _GEN_363,
  output        _GEN_320,
  output        _GEN_314,
  output        _GEN_329,
  output        _GEN_321_0,
  output        _GEN_327_0,
  output        _GEN_103_0,
  output        _GEN_97,
  output        _GEN_236,
  output        _GEN_354,
  output        _GEN_234_0,
  output        _GEN_130,
  output        _GEN_61,
  output        _GEN_55,
  output        _GEN_249_0,
  output        _GEN_335,
  output        _GEN_243,
  output        _GEN_447,
  output        _GEN_158,
  output        _GEN_330_0,
  output        _GEN_422,
  output        _GEN_245,
  output        _GEN_37,
  output        _GEN_125_0,
  output        _GEN_429,
  output        _GEN_70,
  output        _GEN_64,
  output        _GEN_344,
  output        _GEN_338,
  output        _GEN_293_0,
  output        _GEN_87,
  output        _GEN_416,
  output        _GEN_406_0,
  output        _GEN_58,
  output        _GEN_414_0,
  output        _GEN_309,
  output        _GEN_85_0,
  output        _GEN_299_0,
  output        _GEN_336,
  output        _GEN_408,
  output        _GEN_112,
  output        _GEN_43,
  output        _GEN_150,
  output        _GEN_131,
  output        _GEN_435,
  output        _GEN_230,
  output        _GEN_97_0,
  output        _GEN_124,
  output        _GEN_239,
  output        _GEN_118,
  output        _GEN_392_0,
  output        _GEN_398_0,
  output        _GEN_423_0,
  output        _GEN_237,
  output        _GEN_152,
  output        _GEN_307_0,
  output        _GEN_146_0,
  output        _GEN_315_0,
  output        _GEN_79,
  output        _GEN_224,
  output        _GEN_110,
  output        _GEN_119_0,
  output        _GEN_323,
  output        _GEN_317,
  output        _GEN_79_0,
  output        _GEN_218,
  output        _GEN_208,
  output        _GEN_1_1,
  output        _GEN_196,
  output        _GEN_90,
  output        _GEN_31,
  output        _GEN_400,
  output        _GEN_113_0,
  output        _GEN_162,
  output        _GEN_212,
  output        _GEN_302_0,
  output        _GEN_181,
  output        _GEN_106_0,
  output        _GEN_227,
  output        _GEN_71_0,
  output        _GEN_380_0,
  output        _GEN_425,
  output        _GEN_280,
  output        _GEN_46,
  output        _GEN_174,
  output        _GEN_134,
  output        _GEN_289,
  output        _GEN_318_0,
  output        _GEN_287_0,
  output        _GEN_202,
  output        _GEN_419,
  output        _GEN_388,
  output        _GEN_410,
  output        _GEN_386_0,
  output        _GEN_52,
  output        _GEN_311,
  output        _GEN_301,
  output        _GEN_295,
  output        _GEN_67,
  output        _GEN_281_0,
  output        _GEN_312_0,
  output        _GEN_25,
  output        _GEN_409_0,
  output        _GEN_417_0,
  output        _GEN_411_0,
  output        _GEN_326,
  output        _GEN_55_0,
  output        _GEN_100_0,
  output        _GEN_394,
  output        _GEN_168_0,
  output        _GEN_128,
  output        _GEN_401_0,
  output        _GEN_44_0,
  output        _GEN_376,
  output        _GEN_74_0,
  output        _GEN_374_0,
  output        _GEN_40,
  output        _GEN_368_0,
  output        _GEN_34,
  output        _GEN_383_0,
  output        _GEN_49,
  output        _GEN_263_0,
  output        _GEN_177,
  output        _GEN_171,
  output        _GEN_446,
  output        _GEN_102,
  output        _GEN_290_0,
  output        _GEN_190,
  output        _GEN_83,
  output        _GEN_205,
  output        _GEN_135_0,
  output        _GEN_389_0,
  output        _GEN_93,
  output        _GEN_254_0,
  output        _GEN_298,
  output        _GEN_163_0,
  output        _GEN_21,
  output        _GEN_461,
  output        _GEN_362_0,
  output        _GEN_14,
  output        _GEN_116,
  output        _GEN_156,
  output        _GEN_150_0,
  output        _GEN_283,
  output        _GEN_184,
  output        _GEN_178_0,
  output        _GEN_68_0,
  output        _GEN_296_0,
  output        _GEN_382,
  output        _GEN_397,
  output        _GEN_277,
  output        _GEN_395_0,
  output        _GEN_304_0,
  output        _GEN_199,
  output        _GEN_403,
  output        _GEN_262,
  output        _GEN_28,
  output        _GEN_275_0,
  output        _GEN_269_0,
  output        _GEN_361,
  output        _GEN_96,
  output        _GEN_278_0,
  output        _GEN_193,
  output        _GEN_379,
  output        _GEN_244_0,
  output        _GEN_138,
  output        _GEN_271,
  output        _GEN_251_0,
  output        _GEN_151_1,
  output        _GEN_166_0,
  output        _GEN_455,
  output        _GEN_370,
  output        _GEN_364,
  output        _GEN_259,
  output        _GEN_377_0,
  output        _GEN_153_0,
  output        _GEN_292,
  output        _GEN_84,
  output        _GEN_78,
  output        _GEN_272_0,
  output        _GEN_47_0,
  output        _GEN_335_0,
  output        _GEN_41_0,
  output        _GEN_385,
  output        _GEN_250,
  output        _GEN_434,
  output        _GEN_257_0,
  output        _GEN_343,
  output        _GEN_443,
  output        _GEN_105,
  output        _GEN_99,
  output        _GEN_358,
  output        _GEN_356_0,
  output        _GEN_350_0,
  output        _GEN_132_0,
  output        _GEN_22,
  output        _GEN_144,
  output        _GEN_265,
  output        _GEN_17,
  output        _GEN_159,
  output        _GEN_428,
  output        _GEN_449,
  output        _GEN_90_0,
  output        _GEN_172_0,
  output        _GEN_187,
  output        _GEN_117_0,
  output        _GEN_236_0,
  output        _GEN_371_0,
  output        _GEN_391,
  output        _GEN_165,
  output        _GEN_286,
  output        _GEN_145_0,
  output        _GEN_284_0,
  output        _GEN_232,
  output        _GEN_147_0,
  output        _GEN_416_0,
  output        _GEN_274,
  output        _GEN_260_0,
  output        _GEN_175_0,
  output        _GEN_105_0,
  output        _GEN_169_0,
  output        _GEN_338_0,
  output        _GEN_247,
  output        _GEN_133_0,
  output        _GEN_141_0,
  output        _GEN_160_0,
  output        _GEN_346,
  output        _GEN_99_0,
  output        _GEN_344_0,
  output        _GEN_373,
  output        _GEN_424_0,
  output        _GEN_239_0,
  output        _GEN_353_0,
  output        _GEN_268,
  output        _GEN_127_0,
  output        _GEN_8,
  output        _GEN_266_0,
  output        _GEN_331_0,
  output        _GEN_452,
  output        _GEN_93_0,
  output        _GEN_87_0,
  output        _GEN_367,
  output        _GEN_226,
  output        _GEN_120_0,
  output        _GEN_365_0,
  output        _GEN_6,
  output        _GEN_410_0,
  output        _GEN_253_0,
  output        _GEN_152_0,
  output        _GEN_325_0,
  output        _GEN_148_0,
  output        _GEN_437,
  output        _GEN_352_0,
  output        _GEN_332_0,
  output        _GEN_108,
  output        _GEN_126_0,
  output        _GEN_245_0,
  output        _GEN_359_0,
  output        _GEN_431,
  output        _GEN_72_0,
  output        _GEN_66,
  output        _GEN_154_0,
  output        _GEN_458,
  output        _GEN_317_0,
  output        _GEN_326_0,
  output        _GEN_241,
  output        _GEN_341_0,
  output        _GEN_402_0,
  output        _GEN_1_2,
  output        _GEN_48,
  output        _GEN_394_0,
  output        _GEN_60,
  output        _GEN_248_0,
  output        _GEN_75_0,
  output        _GEN_349,
  output        _GEN_214,
  output        _GEN_347_0,
  output        _GEN_412_0,
  output        _GEN_92_0,
  output        _GEN_102_0,
  output        _GEN_256,
  output        _GEN_121_0,
  output        _GEN_425_0,
  output        _GEN_305_0,
  output        _GEN_419_0,
  output        _GEN_81,
  output        _GEN_320_0,
  output        _GEN_108_0,
  output        _GEN_114_0,
  output        _GEN_123_0,
  output        _GEN_413_0,
  output        _GEN_54,
  output        _GEN_136_0,
  output        _GEN_142_0,
  output        _GEN_440,
  output        _GEN_295_0,
  output        _GEN_340,
  output        _GEN_355,
  output        _GEN_235,
  output        _GEN_129_0,
  output        _GEN_404_0,
  output        _GEN_403_0,
  output        _GEN_313_0,
  output        _GEN_242_0,
  output        _GEN_69_0,
  output        _GEN_157_0,
  output        _GEN_220,
  output        _GEN_229,
  output        _GEN_115_0,
  output        _GEN_15_0,
  output        _GEN_334,
  output        _GEN_328,
  output        _GEN_96_0,
  output        _GEN_86_0,
  output        _GEN_36,
  output        _GEN_405_0,
  output        _GEN_415_0,
  output        _GEN_164_0,
  output        _GEN_124_0,
  output        _GEN_322,
  output        _GEN_308_0,
  output        _GEN_337_0,
  output        _GEN_223,
  output        _GEN_217,
  output        _GEN_192,
  output        _GEN_390_0,
  output        _GEN_42_0,
  output        _GEN_149_0,
  output        _GEN_291_0,
  output        _GEN_139_0,
  output        _GEN_329_0,
  output        _GEN_292_0,
  output        _GEN_298_0,
  output        _GEN_207,
  output        _GEN_399_0,
  output        _GEN_421,
  output        _GEN_63,
  output        _GEN_391_0,
  output        _GEN_316_0,
  output        _GEN_306_0,
  output        _GEN_314_0,
  output        _GEN_21_0,
  output        _GEN_323_0,
  output        _GEN_384_0,
  output        _GEN_118_0,
  output        _GEN_376_0,
  output        _GEN_422_0,
  output        _GEN_277_0,
  output        _GEN_57,
  output        _GEN_130_0,
  output        _GEN_46_0,
  output        _GEN_111_0,
  output        _GEN_78_0,
  output        _GEN_238_0,
  output        _GEN_407_0,
  output        _GEN_179_0,
  output        _GEN_397_0,
  output        _GEN_173_0,
  output        _GEN_70_0,
  output        _GEN_379_0,
  output        _GEN_82_0,
  output        _GEN_373_0,
  output        _GEN_45_0,
  output        _GEN_54_0,
  output        _GEN_201,
  output        _GEN_195,
  output        _GEN_364_0,
  output        _GEN_259_0,
  output        _GEN_167_0,
  output        _GEN_309_0,
  output        _GEN_43_0,
  output        _GEN_372_0,
  output        _GEN_19,
  output        _GEN_161_0,
  output        _GEN_51,
  output        _GEN_265_0,
  output        _GEN_294_0,
  output        _GEN_180,
  output        _GEN_189,
  output        _GEN_211,
  output        _GEN_301_0,
  output        _GEN_393_0,
  output        _GEN_387_0,
  output        _GEN_39,
  output        _GEN_146_1,
  output        _GEN_288_0,
  output        _GEN_310_0,
  output        _GEN_300_0,
  output        _GEN_286_0,
  output        _GEN_400_0,
  output        _GEN_319_0,
  output        _GEN_107_0,
  output        _GEN_174_0,
  output        _GEN_89,
  output        _GEN_358_0,
  output        _GEN_30,
  output        _GEN_24,
  output        _GEN_408_0,
  output        _GEN_418_0,
  output        _GEN_273_0,
  output        _GEN_5_0,
  output        _GEN_112_0,
  output        _GEN_385_0,
  output        _GEN_457,
  output        _GEN_311_0,
  output        _GEN_280_0,
  output        _GEN_366_0,
  output        _GEN_360_0,
  output        _GEN_354_0,
  output        _GEN_143_0,
  output        _GEN_367_0,
  output        _GEN_33_0,
  output        _GEN_247_0,
  output        _GEN_276_0,
  output        _GEN_348_0,
  output        _GEN_274_0,
  output        _GEN_460,
  output        _GEN_101_0,
  output        _GEN_375_0,
  output        _GEN_283_0,
  output        _GEN_27,
  output        _GEN_13,
  output        _GEN_388_0,
  output        _GEN_382_0,
  output        _GEN_268_0,
  output        _GEN_297_0,
  output        _GEN_89_0,
  output        _GEN_176_0,
  output        _GEN_177_0,
  output        _GEN_346_0,
  output        _GEN_64_0,
  output        _GEN_340_0,
  output        _GEN_255_0,
  output        _GEN_204,
  output        _GEN_134_0,
  output        _GEN_149_1,
  output        _GEN_439,
  output        _GEN_80_0,
  output        _GEN_262_0,
  output        _GEN_303_0,
  output        _GEN_162_0,
  output        _GEN_17_0,
  output        _GEN_198,
  output        _GEN_361_0,
  output        _GEN_381_0,
  output        _GEN_261_0,
  output        _GEN_155_0,
  output        _GEN_156_0,
  output        _GEN_170_0,
  output        _GEN_95_0,
  output        _GEN_183,
  output        _GEN_369_0,
  output        _GEN_73_0,
  output        _GEN_128_0,
  output        _GEN_241_0,
  output        _GEN_282_0,
  output        _GEN_396_0,
  output        _GEN_445,
  output        _GEN_289_0,
  output        _GEN_378_0,
  output        _GEN_186,
  output        _GEN_131_0,
  output        _GEN_152_1,
  output        _GEN_421_0,
  output        _GEN_427,
  output        _GEN_62,
  output        _GEN_285_0,
  output        _GEN_336_0,
  output        _GEN_144_0,
  output        _GEN_150_1,
  output        _GEN_454,
  output        _GEN_363_0,
  output        _GEN_243_0,
  output        _GEN_258_0,
  output        _GEN_138_0,
  output        _GEN_256_0,
  output        _GEN_171_0,
  output        _GEN_357_0,
  output        _GEN_165_0,
  output        _GEN_110_0,
  output        _GEN_40_0,
  output        _GEN_264_0,
  output        _GEN_5_1,
  output        _GEN_158_0,
  output        _GEN_16_0,
  output        _GEN_271_0,
  output        _GEN_342_0,
  output        _GEN_322_0,
  output        _GEN_98_0,
  output        _GEN_237_0,
  output        _GEN_334_0,
  output        _GEN_116_0,
  output        _GEN_235_0,
  output        _GEN_349_0,
  output        _GEN_147_1,
  output        _GEN_448,
  output        _GEN_442,
  output        _GEN_83_0,
  output        _GEN_343_0,
  output        _GEN_355_0,
  output        _GEN_137_0,
  output        _GEN_370_0,
  output        _GEN_250_0,
  output        _GEN_77,
  output        _GEN_270_0,
  output        _GEN_279_0,
  output        _GEN_159_0,
  output        _GEN_463,
  output        _GEN_328_0,
  output        _GEN_104_0
);
  wire  c_metaReset; // @[core.scala 24:19]
  wire  c_clock; // @[core.scala 24:19]
  wire  c_reset; // @[core.scala 24:19]
  wire  c_io_imem_resp_valid; // @[core.scala 24:19]
  wire  c_io_dmem_resp_valid; // @[core.scala 24:19]
  wire [31:0] c_io_dat_dec_inst; // @[core.scala 24:19]
  wire  c_io_dat_exe_br_eq; // @[core.scala 24:19]
  wire  c_io_dat_exe_br_lt; // @[core.scala 24:19]
  wire  c_io_dat_exe_br_ltu; // @[core.scala 24:19]
  wire [3:0] c_io_dat_exe_br_type; // @[core.scala 24:19]
  wire  c_io_dat_mem_ctrl_dmem_val; // @[core.scala 24:19]
  wire  c_io_dat_csr_eret; // @[core.scala 24:19]
  wire  c_io_ctl_dec_stall; // @[core.scala 24:19]
  wire  c_io_ctl_full_stall; // @[core.scala 24:19]
  wire [1:0] c_io_ctl_exe_pc_sel; // @[core.scala 24:19]
  wire [3:0] c_io_ctl_br_type; // @[core.scala 24:19]
  wire  c_io_ctl_if_kill; // @[core.scala 24:19]
  wire  c_io_ctl_dec_kill; // @[core.scala 24:19]
  wire [1:0] c_io_ctl_op1_sel; // @[core.scala 24:19]
  wire [2:0] c_io_ctl_op2_sel; // @[core.scala 24:19]
  wire [3:0] c_io_ctl_alu_fun; // @[core.scala 24:19]
  wire [1:0] c_io_ctl_wb_sel; // @[core.scala 24:19]
  wire  c_io_ctl_rf_wen; // @[core.scala 24:19]
  wire  c_io_ctl_mem_val; // @[core.scala 24:19]
  wire [1:0] c_io_ctl_mem_fcn; // @[core.scala 24:19]
  wire [2:0] c_io_ctl_mem_typ; // @[core.scala 24:19]
  wire [2:0] c_io_ctl_csr_cmd; // @[core.scala 24:19]
  wire  c_io_ctl_fencei; // @[core.scala 24:19]
  wire  c_io_ctl_pipeline_kill; // @[core.scala 24:19]
  wire  c_io_ctl_mem_exception; // @[core.scala 24:19]
  wire  c__GEN_111_0; // @[core.scala 24:19]
  wire  c__GEN_71_0; // @[core.scala 24:19]
  wire  c__GEN_324_0; // @[core.scala 24:19]
  wire  c__GEN_219_0; // @[core.scala 24:19]
  wire  c__GEN_168_0; // @[core.scala 24:19]
  wire  c__GEN_1_0; // @[core.scala 24:19]
  wire  c__GEN_423_0; // @[core.scala 24:19]
  wire  c__GEN_44_0; // @[core.scala 24:19]
  wire  c__GEN_267_0; // @[core.scala 24:19]
  wire  c__GEN_126_0; // @[core.scala 24:19]
  wire  c__GEN_153_0; // @[core.scala 24:19]
  wire  c__GEN_225_0; // @[core.scala 24:19]
  wire  c__GEN_59_0; // @[core.scala 24:19]
  wire  c__GEN_252_0; // @[core.scala 24:19]
  wire  c__GEN_147_0; // @[core.scala 24:19]
  wire  c__GEN_351_0; // @[core.scala 24:19]
  wire  c__GEN_210_0; // @[core.scala 24:19]
  wire  c__GEN_246_0; // @[core.scala 24:19]
  wire  c__GEN_65_0; // @[core.scala 24:19]
  wire  c__GEN_132_0; // @[core.scala 24:19]
  wire  c__GEN_318_0; // @[core.scala 24:19]
  wire  c__GEN_92_0; // @[core.scala 24:19]
  wire  c__GEN_345_0; // @[core.scala 24:19]
  wire  c__GEN_231_0; // @[core.scala 24:19]
  wire  c__GEN_417_0; // @[core.scala 24:19]
  wire  c__GEN_50_0; // @[core.scala 24:19]
  wire  c__GEN_330_0; // @[core.scala 24:19]
  wire  c__GEN_86_0; // @[core.scala 24:19]
  wire  c__GEN_339_0; // @[core.scala 24:19]
  wire  c__GEN_240_0; // @[core.scala 24:19]
  wire  c__GEN_234_0; // @[core.scala 24:19]
  wire  c__GEN_120_0; // @[core.scala 24:19]
  wire  c__GEN_129_0; // @[core.scala 24:19]
  wire  c__GEN_333_0; // @[core.scala 24:19]
  wire  c__GEN_302_0; // @[core.scala 24:19]
  wire  c__GEN_228_0; // @[core.scala 24:19]
  wire  c__GEN_197_0; // @[core.scala 24:19]
  wire  c__GEN_411_0; // @[core.scala 24:19]
  wire  c__GEN_401_0; // @[core.scala 24:19]
  wire  c__GEN_47_0; // @[core.scala 24:19]
  wire  c__GEN_296_0; // @[core.scala 24:19]
  wire  c__GEN_74_0; // @[core.scala 24:19]
  wire  c__GEN_213_0; // @[core.scala 24:19]
  wire  c__GEN_32_0; // @[core.scala 24:19]
  wire  c__GEN_68_0; // @[core.scala 24:19]
  wire  c__GEN_135_0; // @[core.scala 24:19]
  wire  c__GEN_26_0; // @[core.scala 24:19]
  wire  c__GEN_53_0; // @[core.scala 24:19]
  wire  c__GEN_141_0; // @[core.scala 24:19]
  wire  c__GEN_327_0; // @[core.scala 24:19]
  wire  c__GEN_395_0; // @[core.scala 24:19]
  wire  c__GEN_249_0; // @[core.scala 24:19]
  wire  c__GEN_114_0; // @[core.scala 24:19]
  wire  c__GEN_312_0; // @[core.scala 24:19]
  wire  c__GEN_203_0; // @[core.scala 24:19]
  wire  c__GEN_20_0; // @[core.scala 24:19]
  wire  c__GEN_15_0; // @[core.scala 24:19]
  wire  c__GEN_216_0; // @[core.scala 24:19]
  wire  c__GEN_206_0; // @[core.scala 24:19]
  wire  c__GEN_420_0; // @[core.scala 24:19]
  wire  c__GEN_123_0; // @[core.scala 24:19]
  wire  c__GEN_315_0; // @[core.scala 24:19]
  wire  c__GEN_284_0; // @[core.scala 24:19]
  wire  c__GEN_179_0; // @[core.scala 24:19]
  wire  c__GEN_222_0; // @[core.scala 24:19]
  wire  c__GEN_377_0; // @[core.scala 24:19]
  wire  c__GEN_191_0; // @[core.scala 24:19]
  wire  c__GEN_290_0; // @[core.scala 24:19]
  wire  c__GEN_404_0; // @[core.scala 24:19]
  wire  c__GEN_56_1; // @[core.scala 24:19]
  wire  c__GEN_305_0; // @[core.scala 24:19]
  wire  c__GEN_299_0; // @[core.scala 24:19]
  wire  c__GEN_185_0; // @[core.scala 24:19]
  wire  c__GEN_398_0; // @[core.scala 24:19]
  wire  c__GEN_41_0; // @[core.scala 24:19]
  wire  c__GEN_321_0; // @[core.scala 24:19]
  wire  c__GEN_414_0; // @[core.scala 24:19]
  wire  c__GEN_383_0; // @[core.scala 24:19]
  wire  c__GEN_35_0; // @[core.scala 24:19]
  wire  c__GEN_29_0; // @[core.scala 24:19]
  wire  c__GEN_278_0; // @[core.scala 24:19]
  wire  c__GEN_117_0; // @[core.scala 24:19]
  wire  c__GEN_365_0; // @[core.scala 24:19]
  wire  c__GEN_359_0; // @[core.scala 24:19]
  wire  c__GEN_38_0; // @[core.scala 24:19]
  wire  c__GEN_167_0; // @[core.scala 24:19]
  wire  c__GEN_350_0; // @[core.scala 24:19]
  wire  c__GEN_106_0; // @[core.scala 24:19]
  wire  c__GEN_18_0; // @[core.scala 24:19]
  wire  c__GEN_293_0; // @[core.scala 24:19]
  wire  c__GEN_371_0; // @[core.scala 24:19]
  wire  c__GEN_251_0; // @[core.scala 24:19]
  wire  c__GEN_209_0; // @[core.scala 24:19]
  wire  c__GEN_308_0; // @[core.scala 24:19]
  wire  c__GEN_173_0; // @[core.scala 24:19]
  wire  c__GEN_200_0; // @[core.scala 24:19]
  wire  c__GEN_386_0; // @[core.scala 24:19]
  wire  c__GEN_272_0; // @[core.scala 24:19]
  wire  c__GEN_91_1; // @[core.scala 24:19]
  wire  c__GEN_194_0; // @[core.scala 24:19]
  wire  c__GEN_188_0; // @[core.scala 24:19]
  wire  c__GEN_392_0; // @[core.scala 24:19]
  wire  c__GEN_23_0; // @[core.scala 24:19]
  wire  c__GEN_407_0; // @[core.scala 24:19]
  wire  c__GEN_287_0; // @[core.scala 24:19]
  wire  c__GEN_266_0; // @[core.scala 24:19]
  wire  c__GEN_374_0; // @[core.scala 24:19]
  wire  c__GEN_233_0; // @[core.scala 24:19]
  wire  c__GEN_269_0; // @[core.scala 24:19]
  wire  c__GEN_260_0; // @[core.scala 24:19]
  wire  c__GEN_161_0; // @[core.scala 24:19]
  wire  c__GEN_155_0; // @[core.scala 24:19]
  wire  c__GEN_368_0; // @[core.scala 24:19]
  wire  c__GEN_254_0; // @[core.scala 24:19]
  wire  c__GEN_281_0; // @[core.scala 24:19]
  wire  c__GEN_73_0; // @[core.scala 24:19]
  wire  c__GEN_353_0; // @[core.scala 24:19]
  wire  c__GEN_332_0; // @[core.scala 24:19]
  wire  c__GEN_88_1; // @[core.scala 24:19]
  wire  c__GEN_176_0; // @[core.scala 24:19]
  wire  c__GEN_380_0; // @[core.scala 24:19]
  wire  c__GEN_389_0; // @[core.scala 24:19]
  wire  c__GEN_94_0; // @[core.scala 24:19]
  wire  c__GEN_347_0; // @[core.scala 24:19]
  wire  c__GEN_109_0; // @[core.scala 24:19]
  wire  c__GEN_182_0; // @[core.scala 24:19]
  wire  c__GEN_9_0; // @[core.scala 24:19]
  wire  c__GEN_149_0; // @[core.scala 24:19]
  wire  c__GEN_248_0; // @[core.scala 24:19]
  wire  c__GEN_275_0; // @[core.scala 24:19]
  wire  c__GEN_140_1; // @[core.scala 24:19]
  wire  c__GEN_100_0; // @[core.scala 24:19]
  wire  c__GEN_362_0; // @[core.scala 24:19]
  wire  c__GEN_413_0; // @[core.scala 24:19]
  wire  c__GEN_76_0; // @[core.scala 24:19]
  wire  c__GEN_164_0; // @[core.scala 24:19]
  wire  c__GEN_242_0; // @[core.scala 24:19]
  wire  c__GEN_137_0; // @[core.scala 24:19]
  wire  c__GEN_341_0; // @[core.scala 24:19]
  wire  c__GEN_263_0; // @[core.scala 24:19]
  wire  c__GEN_257_0; // @[core.scala 24:19]
  wire  c__GEN_122_1; // @[core.scala 24:19]
  wire  c__GEN_143_0; // @[core.scala 24:19]
  wire  c__GEN_82_0; // @[core.scala 24:19]
  wire  c__GEN_170_0; // @[core.scala 24:19]
  wire  c__GEN_356_0; // @[core.scala 24:19]
  wire  c__GEN_221_0; // @[core.scala 24:19]
  wire  c__GEN_215_0; // @[core.scala 24:19]
  wire  c__GEN_320_0; // @[core.scala 24:19]
  wire  c__GEN_314_0; // @[core.scala 24:19]
  wire  c__GEN_329_0; // @[core.scala 24:19]
  wire  c__GEN_103_1; // @[core.scala 24:19]
  wire  c__GEN_97_0; // @[core.scala 24:19]
  wire  c__GEN_236_0; // @[core.scala 24:19]
  wire  c__GEN_61_0; // @[core.scala 24:19]
  wire  c__GEN_55_0; // @[core.scala 24:19]
  wire  c__GEN_335_0; // @[core.scala 24:19]
  wire  c__GEN_158_0; // @[core.scala 24:19]
  wire  c__GEN_422_0; // @[core.scala 24:19]
  wire  c__GEN_245_0; // @[core.scala 24:19]
  wire  c__GEN_37_0; // @[core.scala 24:19]
  wire  c__GEN_125_1; // @[core.scala 24:19]
  wire  c__GEN_70_0; // @[core.scala 24:19]
  wire  c__GEN_64_0; // @[core.scala 24:19]
  wire  c__GEN_344_0; // @[core.scala 24:19]
  wire  c__GEN_338_0; // @[core.scala 24:19]
  wire  c__GEN_416_0; // @[core.scala 24:19]
  wire  c__GEN_406_1; // @[core.scala 24:19]
  wire  c__GEN_58_0; // @[core.scala 24:19]
  wire  c__GEN_85_1; // @[core.scala 24:19]
  wire  c__GEN_43_0; // @[core.scala 24:19]
  wire  c__GEN_131_0; // @[core.scala 24:19]
  wire  c__GEN_230_0; // @[core.scala 24:19]
  wire  c__GEN_239_0; // @[core.scala 24:19]
  wire  c__GEN_152_0; // @[core.scala 24:19]
  wire  c__GEN_307_1; // @[core.scala 24:19]
  wire  c__GEN_146_1; // @[core.scala 24:19]
  wire  c__GEN_224_0; // @[core.scala 24:19]
  wire  c__GEN_110_0; // @[core.scala 24:19]
  wire  c__GEN_119_1; // @[core.scala 24:19]
  wire  c__GEN_323_0; // @[core.scala 24:19]
  wire  c__GEN_317_0; // @[core.scala 24:19]
  wire  c__GEN_79_1; // @[core.scala 24:19]
  wire  c__GEN_218_0; // @[core.scala 24:19]
  wire  c__GEN_208_0; // @[core.scala 24:19]
  wire  c__GEN_196_0; // @[core.scala 24:19]
  wire  c__GEN_31_0; // @[core.scala 24:19]
  wire  c__GEN_400_0; // @[core.scala 24:19]
  wire  c__GEN_113_1; // @[core.scala 24:19]
  wire  c__GEN_212_0; // @[core.scala 24:19]
  wire  c__GEN_181_0; // @[core.scala 24:19]
  wire  c__GEN_227_0; // @[core.scala 24:19]
  wire  c__GEN_425_0; // @[core.scala 24:19]
  wire  c__GEN_280_0; // @[core.scala 24:19]
  wire  c__GEN_46_0; // @[core.scala 24:19]
  wire  c__GEN_134_0; // @[core.scala 24:19]
  wire  c__GEN_289_0; // @[core.scala 24:19]
  wire  c__GEN_202_0; // @[core.scala 24:19]
  wire  c__GEN_419_0; // @[core.scala 24:19]
  wire  c__GEN_388_0; // @[core.scala 24:19]
  wire  c__GEN_410_0; // @[core.scala 24:19]
  wire  c__GEN_52_0; // @[core.scala 24:19]
  wire  c__GEN_311_0; // @[core.scala 24:19]
  wire  c__GEN_301_0; // @[core.scala 24:19]
  wire  c__GEN_295_0; // @[core.scala 24:19]
  wire  c__GEN_67_0; // @[core.scala 24:19]
  wire  c__GEN_25_0; // @[core.scala 24:19]
  wire  c__GEN_409_1; // @[core.scala 24:19]
  wire  c__GEN_326_0; // @[core.scala 24:19]
  wire  c__GEN_394_0; // @[core.scala 24:19]
  wire  c__GEN_128_0; // @[core.scala 24:19]
  wire  c__GEN_376_0; // @[core.scala 24:19]
  wire  c__GEN_40_0; // @[core.scala 24:19]
  wire  c__GEN_34_0; // @[core.scala 24:19]
  wire  c__GEN_49_0; // @[core.scala 24:19]
  wire  c__GEN_102_0; // @[core.scala 24:19]
  wire  c__GEN_190_0; // @[core.scala 24:19]
  wire  c__GEN_205_0; // @[core.scala 24:19]
  wire  c__GEN_298_0; // @[core.scala 24:19]
  wire  c__GEN_163_1; // @[core.scala 24:19]
  wire  c__GEN_14_0; // @[core.scala 24:19]
  wire  c__GEN_116_0; // @[core.scala 24:19]
  wire  c__GEN_283_0; // @[core.scala 24:19]
  wire  c__GEN_184_0; // @[core.scala 24:19]
  wire  c__GEN_178_1; // @[core.scala 24:19]
  wire  c__GEN_382_0; // @[core.scala 24:19]
  wire  c__GEN_397_0; // @[core.scala 24:19]
  wire  c__GEN_277_0; // @[core.scala 24:19]
  wire  c__GEN_304_1; // @[core.scala 24:19]
  wire  c__GEN_199_0; // @[core.scala 24:19]
  wire  c__GEN_403_0; // @[core.scala 24:19]
  wire  c__GEN_262_0; // @[core.scala 24:19]
  wire  c__GEN_28_0; // @[core.scala 24:19]
  wire  c__GEN_361_0; // @[core.scala 24:19]
  wire  c__GEN_96_0; // @[core.scala 24:19]
  wire  c__GEN_193_0; // @[core.scala 24:19]
  wire  c__GEN_379_0; // @[core.scala 24:19]
  wire  c__GEN_244_1; // @[core.scala 24:19]
  wire  c__GEN_271_0; // @[core.scala 24:19]
  wire  c__GEN_151_2; // @[core.scala 24:19]
  wire  c__GEN_166_1; // @[core.scala 24:19]
  wire  c__GEN_370_0; // @[core.scala 24:19]
  wire  c__GEN_364_0; // @[core.scala 24:19]
  wire  c__GEN_259_0; // @[core.scala 24:19]
  wire  c__GEN_292_0; // @[core.scala 24:19]
  wire  c__GEN_84_0; // @[core.scala 24:19]
  wire  c__GEN_78_0; // @[core.scala 24:19]
  wire  c__GEN_385_0; // @[core.scala 24:19]
  wire  c__GEN_250_0; // @[core.scala 24:19]
  wire  c__GEN_343_0; // @[core.scala 24:19]
  wire  c__GEN_105_0; // @[core.scala 24:19]
  wire  c__GEN_99_0; // @[core.scala 24:19]
  wire  c__GEN_358_0; // @[core.scala 24:19]
  wire  c__GEN_22_0; // @[core.scala 24:19]
  wire  c__GEN_265_0; // @[core.scala 24:19]
  wire  c__GEN_17_0; // @[core.scala 24:19]
  wire  c__GEN_90_1; // @[core.scala 24:19]
  wire  c__GEN_172_1; // @[core.scala 24:19]
  wire  c__GEN_187_0; // @[core.scala 24:19]
  wire  c__GEN_391_0; // @[core.scala 24:19]
  wire  c__GEN_286_0; // @[core.scala 24:19]
  wire  c__GEN_145_1; // @[core.scala 24:19]
  wire  c__GEN_232_0; // @[core.scala 24:19]
  wire  c__GEN_274_0; // @[core.scala 24:19]
  wire  c__GEN_175_1; // @[core.scala 24:19]
  wire  c__GEN_169_1; // @[core.scala 24:19]
  wire  c__GEN_247_0; // @[core.scala 24:19]
  wire  c__GEN_133_1; // @[core.scala 24:19]
  wire  c__GEN_160_1; // @[core.scala 24:19]
  wire  c__GEN_346_0; // @[core.scala 24:19]
  wire  c__GEN_373_0; // @[core.scala 24:19]
  wire  c__GEN_424_1; // @[core.scala 24:19]
  wire  c__GEN_268_0; // @[core.scala 24:19]
  wire  c__GEN_127_1; // @[core.scala 24:19]
  wire  c__GEN_8_0; // @[core.scala 24:19]
  wire  c__GEN_331_1; // @[core.scala 24:19]
  wire  c__GEN_93_1; // @[core.scala 24:19]
  wire  c__GEN_87_1; // @[core.scala 24:19]
  wire  c__GEN_367_0; // @[core.scala 24:19]
  wire  c__GEN_226_0; // @[core.scala 24:19]
  wire  c__GEN_253_1; // @[core.scala 24:19]
  wire  c__GEN_325_1; // @[core.scala 24:19]
  wire  c__GEN_148_1; // @[core.scala 24:19]
  wire  c__GEN_352_1; // @[core.scala 24:19]
  wire  c__GEN_108_0; // @[core.scala 24:19]
  wire  c__GEN_72_1; // @[core.scala 24:19]
  wire  c__GEN_66_0; // @[core.scala 24:19]
  wire  c__GEN_154_1; // @[core.scala 24:19]
  wire  c__GEN_241_0; // @[core.scala 24:19]
  wire  c__GEN_402_1; // @[core.scala 24:19]
  wire  c__GEN_48_0; // @[core.scala 24:19]
  wire  c__GEN_60_0; // @[core.scala 24:19]
  wire  c__GEN_75_1; // @[core.scala 24:19]
  wire  c__GEN_349_0; // @[core.scala 24:19]
  wire  c__GEN_214_0; // @[core.scala 24:19]
  wire  c__GEN_412_1; // @[core.scala 24:19]
  wire  c__GEN_256_0; // @[core.scala 24:19]
  wire  c__GEN_121_1; // @[core.scala 24:19]
  wire  c__GEN_81_0; // @[core.scala 24:19]
  wire  c__GEN_54_0; // @[core.scala 24:19]
  wire  c__GEN_136_1; // @[core.scala 24:19]
  wire  c__GEN_142_1; // @[core.scala 24:19]
  wire  c__GEN_340_0; // @[core.scala 24:19]
  wire  c__GEN_355_0; // @[core.scala 24:19]
  wire  c__GEN_235_0; // @[core.scala 24:19]
  wire  c__GEN_313_1; // @[core.scala 24:19]
  wire  c__GEN_69_1; // @[core.scala 24:19]
  wire  c__GEN_157_1; // @[core.scala 24:19]
  wire  c__GEN_220_0; // @[core.scala 24:19]
  wire  c__GEN_229_0; // @[core.scala 24:19]
  wire  c__GEN_115_1; // @[core.scala 24:19]
  wire  c__GEN_334_0; // @[core.scala 24:19]
  wire  c__GEN_328_0; // @[core.scala 24:19]
  wire  c__GEN_36_0; // @[core.scala 24:19]
  wire  c__GEN_405_1; // @[core.scala 24:19]
  wire  c__GEN_415_1; // @[core.scala 24:19]
  wire  c__GEN_124_1; // @[core.scala 24:19]
  wire  c__GEN_322_0; // @[core.scala 24:19]
  wire  c__GEN_337_1; // @[core.scala 24:19]
  wire  c__GEN_223_0; // @[core.scala 24:19]
  wire  c__GEN_217_0; // @[core.scala 24:19]
  wire  c__GEN_192_0; // @[core.scala 24:19]
  wire  c__GEN_390_1; // @[core.scala 24:19]
  wire  c__GEN_42_1; // @[core.scala 24:19]
  wire  c__GEN_291_1; // @[core.scala 24:19]
  wire  c__GEN_139_1; // @[core.scala 24:19]
  wire  c__GEN_207_0; // @[core.scala 24:19]
  wire  c__GEN_399_1; // @[core.scala 24:19]
  wire  c__GEN_421_0; // @[core.scala 24:19]
  wire  c__GEN_63_0; // @[core.scala 24:19]
  wire  c__GEN_316_1; // @[core.scala 24:19]
  wire  c__GEN_306_1; // @[core.scala 24:19]
  wire  c__GEN_21_1; // @[core.scala 24:19]
  wire  c__GEN_384_1; // @[core.scala 24:19]
  wire  c__GEN_118_1; // @[core.scala 24:19]
  wire  c__GEN_57_0; // @[core.scala 24:19]
  wire  c__GEN_130_1; // @[core.scala 24:19]
  wire  c__GEN_238_1; // @[core.scala 24:19]
  wire  c__GEN_45_1; // @[core.scala 24:19]
  wire  c__GEN_201_0; // @[core.scala 24:19]
  wire  c__GEN_195_0; // @[core.scala 24:19]
  wire  c__GEN_309_1; // @[core.scala 24:19]
  wire  c__GEN_372_1; // @[core.scala 24:19]
  wire  c__GEN_19_0; // @[core.scala 24:19]
  wire  c__GEN_51_0; // @[core.scala 24:19]
  wire  c__GEN_294_1; // @[core.scala 24:19]
  wire  c__GEN_180_0; // @[core.scala 24:19]
  wire  c__GEN_189_0; // @[core.scala 24:19]
  wire  c__GEN_211_0; // @[core.scala 24:19]
  wire  c__GEN_393_1; // @[core.scala 24:19]
  wire  c__GEN_387_1; // @[core.scala 24:19]
  wire  c__GEN_39_0; // @[core.scala 24:19]
  wire  c__GEN_288_1; // @[core.scala 24:19]
  wire  c__GEN_310_1; // @[core.scala 24:19]
  wire  c__GEN_300_1; // @[core.scala 24:19]
  wire  c__GEN_319_1; // @[core.scala 24:19]
  wire  c__GEN_107_1; // @[core.scala 24:19]
  wire  c__GEN_174_1; // @[core.scala 24:19]
  wire  c__GEN_30_0; // @[core.scala 24:19]
  wire  c__GEN_24_0; // @[core.scala 24:19]
  wire  c__GEN_408_1; // @[core.scala 24:19]
  wire  c__GEN_418_1; // @[core.scala 24:19]
  wire  c__GEN_273_1; // @[core.scala 24:19]
  wire  c__GEN_5_1; // @[core.scala 24:19]
  wire  c__GEN_112_1; // @[core.scala 24:19]
  wire  c__GEN_366_1; // @[core.scala 24:19]
  wire  c__GEN_360_1; // @[core.scala 24:19]
  wire  c__GEN_354_1; // @[core.scala 24:19]
  wire  c__GEN_33_1; // @[core.scala 24:19]
  wire  c__GEN_276_1; // @[core.scala 24:19]
  wire  c__GEN_348_1; // @[core.scala 24:19]
  wire  c__GEN_101_1; // @[core.scala 24:19]
  wire  c__GEN_375_1; // @[core.scala 24:19]
  wire  c__GEN_27_0; // @[core.scala 24:19]
  wire  c__GEN_13_0; // @[core.scala 24:19]
  wire  c__GEN_297_1; // @[core.scala 24:19]
  wire  c__GEN_89_1; // @[core.scala 24:19]
  wire  c__GEN_177_1; // @[core.scala 24:19]
  wire  c__GEN_255_1; // @[core.scala 24:19]
  wire  c__GEN_204_0; // @[core.scala 24:19]
  wire  c__GEN_80_1; // @[core.scala 24:19]
  wire  c__GEN_303_1; // @[core.scala 24:19]
  wire  c__GEN_162_1; // @[core.scala 24:19]
  wire  c__GEN_198_0; // @[core.scala 24:19]
  wire  c__GEN_381_1; // @[core.scala 24:19]
  wire  c__GEN_261_1; // @[core.scala 24:19]
  wire  c__GEN_156_1; // @[core.scala 24:19]
  wire  c__GEN_95_1; // @[core.scala 24:19]
  wire  c__GEN_183_0; // @[core.scala 24:19]
  wire  c__GEN_369_1; // @[core.scala 24:19]
  wire  c__GEN_282_1; // @[core.scala 24:19]
  wire  c__GEN_396_1; // @[core.scala 24:19]
  wire  c__GEN_378_1; // @[core.scala 24:19]
  wire  c__GEN_186_0; // @[core.scala 24:19]
  wire  c__GEN_62_0; // @[core.scala 24:19]
  wire  c__GEN_285_1; // @[core.scala 24:19]
  wire  c__GEN_336_1; // @[core.scala 24:19]
  wire  c__GEN_144_1; // @[core.scala 24:19]
  wire  c__GEN_150_2; // @[core.scala 24:19]
  wire  c__GEN_363_1; // @[core.scala 24:19]
  wire  c__GEN_243_1; // @[core.scala 24:19]
  wire  c__GEN_258_1; // @[core.scala 24:19]
  wire  c__GEN_138_1; // @[core.scala 24:19]
  wire  c__GEN_171_1; // @[core.scala 24:19]
  wire  c__GEN_357_1; // @[core.scala 24:19]
  wire  c__GEN_165_1; // @[core.scala 24:19]
  wire  c__GEN_264_1; // @[core.scala 24:19]
  wire  c__GEN_16_1; // @[core.scala 24:19]
  wire  c__GEN_342_1; // @[core.scala 24:19]
  wire  c__GEN_98_1; // @[core.scala 24:19]
  wire  c__GEN_237_1; // @[core.scala 24:19]
  wire  c__GEN_83_1; // @[core.scala 24:19]
  wire  c__GEN_77_0; // @[core.scala 24:19]
  wire  c__GEN_270_1; // @[core.scala 24:19]
  wire  c__GEN_279_1; // @[core.scala 24:19]
  wire  c__GEN_159_1; // @[core.scala 24:19]
  wire  c__GEN_104_1; // @[core.scala 24:19]
  wire  d_metaReset; // @[core.scala 25:19]
  wire  d_clock; // @[core.scala 25:19]
  wire  d_reset; // @[core.scala 25:19]
  wire [31:0] d_io_imem_req_bits_addr; // @[core.scala 25:19]
  wire [31:0] d_io_imem_resp_bits_data; // @[core.scala 25:19]
  wire  d_io_dmem_req_valid; // @[core.scala 25:19]
  wire [31:0] d_io_dmem_req_bits_addr; // @[core.scala 25:19]
  wire [31:0] d_io_dmem_req_bits_data; // @[core.scala 25:19]
  wire  d_io_dmem_req_bits_fcn; // @[core.scala 25:19]
  wire [2:0] d_io_dmem_req_bits_typ; // @[core.scala 25:19]
  wire [31:0] d_io_dmem_resp_bits_data; // @[core.scala 25:19]
  wire  d_io_ctl_dec_stall; // @[core.scala 25:19]
  wire  d_io_ctl_full_stall; // @[core.scala 25:19]
  wire [1:0] d_io_ctl_exe_pc_sel; // @[core.scala 25:19]
  wire [3:0] d_io_ctl_br_type; // @[core.scala 25:19]
  wire  d_io_ctl_if_kill; // @[core.scala 25:19]
  wire  d_io_ctl_dec_kill; // @[core.scala 25:19]
  wire [1:0] d_io_ctl_op1_sel; // @[core.scala 25:19]
  wire [2:0] d_io_ctl_op2_sel; // @[core.scala 25:19]
  wire [3:0] d_io_ctl_alu_fun; // @[core.scala 25:19]
  wire [1:0] d_io_ctl_wb_sel; // @[core.scala 25:19]
  wire  d_io_ctl_rf_wen; // @[core.scala 25:19]
  wire  d_io_ctl_mem_val; // @[core.scala 25:19]
  wire [1:0] d_io_ctl_mem_fcn; // @[core.scala 25:19]
  wire [2:0] d_io_ctl_mem_typ; // @[core.scala 25:19]
  wire [2:0] d_io_ctl_csr_cmd; // @[core.scala 25:19]
  wire  d_io_ctl_fencei; // @[core.scala 25:19]
  wire  d_io_ctl_pipeline_kill; // @[core.scala 25:19]
  wire  d_io_ctl_mem_exception; // @[core.scala 25:19]
  wire [31:0] d_io_dat_dec_inst; // @[core.scala 25:19]
  wire  d_io_dat_exe_br_eq; // @[core.scala 25:19]
  wire  d_io_dat_exe_br_lt; // @[core.scala 25:19]
  wire  d_io_dat_exe_br_ltu; // @[core.scala 25:19]
  wire [3:0] d_io_dat_exe_br_type; // @[core.scala 25:19]
  wire  d_io_dat_mem_ctrl_dmem_val; // @[core.scala 25:19]
  wire  d_io_dat_csr_eret; // @[core.scala 25:19]
  wire  d__GEN_451; // @[core.scala 25:19]
  wire  d__GEN_331; // @[core.scala 25:19]
  wire  d__GEN_337; // @[core.scala 25:19]
  wire  d__GEN_113_0; // @[core.scala 25:19]
  wire  d__GEN_415; // @[core.scala 25:19]
  wire  d__GEN_436; // @[core.scala 25:19]
  wire  d__GEN_140_0; // @[core.scala 25:19]
  wire  d__GEN_98_0; // @[core.scala 25:19]
  wire  d__GEN_352; // @[core.scala 25:19]
  wire  d__GEN_125_0; // @[core.scala 25:19]
  wire  d__GEN_430; // @[core.scala 25:19]
  wire  d__GEN_119_0; // @[core.scala 25:19]
  wire  d__GEN_88_0; // @[core.scala 25:19]
  wire  d__GEN_151_0; // @[core.scala 25:19]
  wire  d__GEN_310; // @[core.scala 25:19]
  wire  d__GEN_104_0; // @[core.scala 25:19]
  wire  d__GEN_409; // @[core.scala 25:19]
  wire  d__GEN_253; // @[core.scala 25:19]
  wire  d__GEN_316; // @[core.scala 25:19]
  wire  d__GEN_244; // @[core.scala 25:19]
  wire  d__GEN_238; // @[core.scala 25:19]
  wire  d__GEN_101_0; // @[core.scala 25:19]
  wire  d__GEN_325; // @[core.scala 25:19]
  wire  d__GEN_169_0; // @[core.scala 25:19]
  wire  d__GEN_433; // @[core.scala 25:19]
  wire  d__GEN_313; // @[core.scala 25:19]
  wire  d__GEN_91_0; // @[core.scala 25:19]
  wire  d__GEN_11_0; // @[core.scala 25:19]
  wire  d__GEN_304; // @[core.scala 25:19]
  wire  d__GEN_294; // @[core.scala 25:19]
  wire  d__GEN_303; // @[core.scala 25:19]
  wire  d__GEN_107_0; // @[core.scala 25:19]
  wire  d__GEN_0_0; // @[core.scala 25:19]
  wire  d__GEN_402; // @[core.scala 25:19]
  wire  d__GEN_412; // @[core.scala 25:19]
  wire  d__GEN_424; // @[core.scala 25:19]
  wire  d__GEN_175_0; // @[core.scala 25:19]
  wire  d__GEN_319; // @[core.scala 25:19]
  wire  d__GEN_288; // @[core.scala 25:19]
  wire  d__GEN_56_0; // @[core.scala 25:19]
  wire  d__GEN_418; // @[core.scala 25:19]
  wire  d__GEN_122_0; // @[core.scala 25:19]
  wire  d__GEN_387; // @[core.scala 25:19]
  wire  d__GEN_72_0; // @[core.scala 25:19]
  wire  d__GEN_75_0; // @[core.scala 25:19]
  wire  d__GEN_85_0; // @[core.scala 25:19]
  wire  d__GEN_178_0; // @[core.scala 25:19]
  wire  d__GEN_157_0; // @[core.scala 25:19]
  wire  d__GEN_462; // @[core.scala 25:19]
  wire  d__GEN_69_0; // @[core.scala 25:19]
  wire  d__GEN_375; // @[core.scala 25:19]
  wire  d__GEN_151_1; // @[core.scala 25:19]
  wire  d__GEN_33_0; // @[core.scala 25:19]
  wire  d__GEN_390; // @[core.scala 25:19]
  wire  d__GEN_307; // @[core.scala 25:19]
  wire  d__GEN_297; // @[core.scala 25:19]
  wire  d__GEN_406; // @[core.scala 25:19]
  wire  d__GEN_270; // @[core.scala 25:19]
  wire  d__GEN_95_0; // @[core.scala 25:19]
  wire  d__GEN_45_0; // @[core.scala 25:19]
  wire  d__GEN_369; // @[core.scala 25:19]
  wire  d__GEN_396; // @[core.scala 25:19]
  wire  d__GEN_172_0; // @[core.scala 25:19]
  wire  d__GEN_276; // @[core.scala 25:19]
  wire  d__GEN_291; // @[core.scala 25:19]
  wire  d__GEN_258; // @[core.scala 25:19]
  wire  d__GEN_372; // @[core.scala 25:19]
  wire  d__GEN_252_0; // @[core.scala 25:19]
  wire  d__GEN_166_0; // @[core.scala 25:19]
  wire  d__GEN_285; // @[core.scala 25:19]
  wire  d__GEN_42_0; // @[core.scala 25:19]
  wire  d__GEN_384; // @[core.scala 25:19]
  wire  d__GEN_378; // @[core.scala 25:19]
  wire  d__GEN_393; // @[core.scala 25:19]
  wire  d__GEN_273; // @[core.scala 25:19]
  wire  d__GEN_456; // @[core.scala 25:19]
  wire  d__GEN_80_0; // @[core.scala 25:19]
  wire  d__GEN_351_0; // @[core.scala 25:19]
  wire  d__GEN_139_0; // @[core.scala 25:19]
  wire  d__GEN_145_0; // @[core.scala 25:19]
  wire  d__GEN_450; // @[core.scala 25:19]
  wire  d__GEN_53_1; // @[core.scala 25:19]
  wire  d__GEN_357; // @[core.scala 25:19]
  wire  d__GEN_160_0; // @[core.scala 25:19]
  wire  d__GEN_279; // @[core.scala 25:19]
  wire  d__GEN_133_0; // @[core.scala 25:19]
  wire  d__GEN_399; // @[core.scala 25:19]
  wire  d__GEN_264; // @[core.scala 25:19]
  wire  d__GEN_300; // @[core.scala 25:19]
  wire  d__GEN_127_0; // @[core.scala 25:19]
  wire  d__GEN_432; // @[core.scala 25:19]
  wire  d__GEN_381; // @[core.scala 25:19]
  wire  d__GEN_339_0; // @[core.scala 25:19]
  wire  d__GEN_261; // @[core.scala 25:19]
  wire  d__GEN_16_0; // @[core.scala 25:19]
  wire  d__GEN_360; // @[core.scala 25:19]
  wire  d__GEN_163_0; // @[core.scala 25:19]
  wire  d__GEN_246_0; // @[core.scala 25:19]
  wire  d__GEN_438; // @[core.scala 25:19]
  wire  d__GEN_282; // @[core.scala 25:19]
  wire  d__GEN_345_0; // @[core.scala 25:19]
  wire  d__GEN_121_0; // @[core.scala 25:19]
  wire  d__GEN_240_0; // @[core.scala 25:19]
  wire  d__GEN_148_0; // @[core.scala 25:19]
  wire  d__GEN_154_0; // @[core.scala 25:19]
  wire  d__GEN_444; // @[core.scala 25:19]
  wire  d__GEN_267_0; // @[core.scala 25:19]
  wire  d__GEN_459; // @[core.scala 25:19]
  wire  d__GEN_453; // @[core.scala 25:19]
  wire  d__GEN_366; // @[core.scala 25:19]
  wire  d__GEN_7_0; // @[core.scala 25:19]
  wire  d__GEN_142_0; // @[core.scala 25:19]
  wire  d__GEN_324_0; // @[core.scala 25:19]
  wire  d__GEN_333_0; // @[core.scala 25:19]
  wire  d__GEN_342; // @[core.scala 25:19]
  wire  d__GEN_405; // @[core.scala 25:19]
  wire  d__GEN_420_0; // @[core.scala 25:19]
  wire  d__GEN_306; // @[core.scala 25:19]
  wire  d__GEN_109_1; // @[core.scala 25:19]
  wire  d__GEN_103_0; // @[core.scala 25:19]
  wire  d__GEN_3_0; // @[core.scala 25:19]
  wire  d__GEN_136_0; // @[core.scala 25:19]
  wire  d__GEN_426; // @[core.scala 25:19]
  wire  d__GEN_441; // @[core.scala 25:19]
  wire  d__GEN_94_1; // @[core.scala 25:19]
  wire  d__GEN_348; // @[core.scala 25:19]
  wire  d__GEN_255; // @[core.scala 25:19]
  wire  d__GEN_115_0; // @[core.scala 25:19]
  wire  d__GEN_146_0; // @[core.scala 25:19]
  wire  d__GEN_363; // @[core.scala 25:19]
  wire  d__GEN_321_0; // @[core.scala 25:19]
  wire  d__GEN_327_0; // @[core.scala 25:19]
  wire  d__GEN_354; // @[core.scala 25:19]
  wire  d__GEN_234_0; // @[core.scala 25:19]
  wire  d__GEN_130_0; // @[core.scala 25:19]
  wire  d__GEN_249_0; // @[core.scala 25:19]
  wire  d__GEN_243; // @[core.scala 25:19]
  wire  d__GEN_447; // @[core.scala 25:19]
  wire  d__GEN_330_0; // @[core.scala 25:19]
  wire  d__GEN_429; // @[core.scala 25:19]
  wire  d__GEN_293_0; // @[core.scala 25:19]
  wire  d__GEN_87_0; // @[core.scala 25:19]
  wire  d__GEN_414_0; // @[core.scala 25:19]
  wire  d__GEN_309; // @[core.scala 25:19]
  wire  d__GEN_299_0; // @[core.scala 25:19]
  wire  d__GEN_336; // @[core.scala 25:19]
  wire  d__GEN_408; // @[core.scala 25:19]
  wire  d__GEN_112_0; // @[core.scala 25:19]
  wire  d__GEN_150_0; // @[core.scala 25:19]
  wire  d__GEN_435; // @[core.scala 25:19]
  wire  d__GEN_97_1; // @[core.scala 25:19]
  wire  d__GEN_124_0; // @[core.scala 25:19]
  wire  d__GEN_118_0; // @[core.scala 25:19]
  wire  d__GEN_392_0; // @[core.scala 25:19]
  wire  d__GEN_398_0; // @[core.scala 25:19]
  wire  d__GEN_423_0; // @[core.scala 25:19]
  wire  d__GEN_237; // @[core.scala 25:19]
  wire  d__GEN_315_0; // @[core.scala 25:19]
  wire  d__GEN_79_0; // @[core.scala 25:19]
  wire  d__GEN_1_2; // @[core.scala 25:19]
  wire  d__GEN_90_0; // @[core.scala 25:19]
  wire  d__GEN_162_0; // @[core.scala 25:19]
  wire  d__GEN_302_0; // @[core.scala 25:19]
  wire  d__GEN_106_1; // @[core.scala 25:19]
  wire  d__GEN_71_1; // @[core.scala 25:19]
  wire  d__GEN_380_0; // @[core.scala 25:19]
  wire  d__GEN_174_0; // @[core.scala 25:19]
  wire  d__GEN_318_0; // @[core.scala 25:19]
  wire  d__GEN_287_0; // @[core.scala 25:19]
  wire  d__GEN_386_0; // @[core.scala 25:19]
  wire  d__GEN_281_0; // @[core.scala 25:19]
  wire  d__GEN_312_0; // @[core.scala 25:19]
  wire  d__GEN_417_0; // @[core.scala 25:19]
  wire  d__GEN_411_0; // @[core.scala 25:19]
  wire  d__GEN_55_1; // @[core.scala 25:19]
  wire  d__GEN_100_1; // @[core.scala 25:19]
  wire  d__GEN_168_1; // @[core.scala 25:19]
  wire  d__GEN_401_0; // @[core.scala 25:19]
  wire  d__GEN_44_1; // @[core.scala 25:19]
  wire  d__GEN_74_1; // @[core.scala 25:19]
  wire  d__GEN_374_0; // @[core.scala 25:19]
  wire  d__GEN_368_0; // @[core.scala 25:19]
  wire  d__GEN_383_0; // @[core.scala 25:19]
  wire  d__GEN_263_0; // @[core.scala 25:19]
  wire  d__GEN_177_0; // @[core.scala 25:19]
  wire  d__GEN_171_0; // @[core.scala 25:19]
  wire  d__GEN_446; // @[core.scala 25:19]
  wire  d__GEN_290_0; // @[core.scala 25:19]
  wire  d__GEN_83_0; // @[core.scala 25:19]
  wire  d__GEN_135_1; // @[core.scala 25:19]
  wire  d__GEN_389_0; // @[core.scala 25:19]
  wire  d__GEN_93_0; // @[core.scala 25:19]
  wire  d__GEN_254_0; // @[core.scala 25:19]
  wire  d__GEN_21_0; // @[core.scala 25:19]
  wire  d__GEN_461; // @[core.scala 25:19]
  wire  d__GEN_362_0; // @[core.scala 25:19]
  wire  d__GEN_156_0; // @[core.scala 25:19]
  wire  d__GEN_150_1; // @[core.scala 25:19]
  wire  d__GEN_68_1; // @[core.scala 25:19]
  wire  d__GEN_296_0; // @[core.scala 25:19]
  wire  d__GEN_395_0; // @[core.scala 25:19]
  wire  d__GEN_275_0; // @[core.scala 25:19]
  wire  d__GEN_269_0; // @[core.scala 25:19]
  wire  d__GEN_278_0; // @[core.scala 25:19]
  wire  d__GEN_138_0; // @[core.scala 25:19]
  wire  d__GEN_251_0; // @[core.scala 25:19]
  wire  d__GEN_455; // @[core.scala 25:19]
  wire  d__GEN_377_0; // @[core.scala 25:19]
  wire  d__GEN_153_1; // @[core.scala 25:19]
  wire  d__GEN_272_0; // @[core.scala 25:19]
  wire  d__GEN_47_1; // @[core.scala 25:19]
  wire  d__GEN_335_0; // @[core.scala 25:19]
  wire  d__GEN_41_1; // @[core.scala 25:19]
  wire  d__GEN_434; // @[core.scala 25:19]
  wire  d__GEN_257_0; // @[core.scala 25:19]
  wire  d__GEN_443; // @[core.scala 25:19]
  wire  d__GEN_356_0; // @[core.scala 25:19]
  wire  d__GEN_350_0; // @[core.scala 25:19]
  wire  d__GEN_132_1; // @[core.scala 25:19]
  wire  d__GEN_144_0; // @[core.scala 25:19]
  wire  d__GEN_159_0; // @[core.scala 25:19]
  wire  d__GEN_428; // @[core.scala 25:19]
  wire  d__GEN_449; // @[core.scala 25:19]
  wire  d__GEN_117_1; // @[core.scala 25:19]
  wire  d__GEN_236_0; // @[core.scala 25:19]
  wire  d__GEN_371_0; // @[core.scala 25:19]
  wire  d__GEN_165_0; // @[core.scala 25:19]
  wire  d__GEN_284_0; // @[core.scala 25:19]
  wire  d__GEN_147_1; // @[core.scala 25:19]
  wire  d__GEN_416_0; // @[core.scala 25:19]
  wire  d__GEN_260_0; // @[core.scala 25:19]
  wire  d__GEN_105_1; // @[core.scala 25:19]
  wire  d__GEN_338_0; // @[core.scala 25:19]
  wire  d__GEN_141_1; // @[core.scala 25:19]
  wire  d__GEN_99_1; // @[core.scala 25:19]
  wire  d__GEN_344_0; // @[core.scala 25:19]
  wire  d__GEN_239_0; // @[core.scala 25:19]
  wire  d__GEN_353_0; // @[core.scala 25:19]
  wire  d__GEN_266_0; // @[core.scala 25:19]
  wire  d__GEN_452; // @[core.scala 25:19]
  wire  d__GEN_120_1; // @[core.scala 25:19]
  wire  d__GEN_365_0; // @[core.scala 25:19]
  wire  d__GEN_6_0; // @[core.scala 25:19]
  wire  d__GEN_410_0; // @[core.scala 25:19]
  wire  d__GEN_152_1; // @[core.scala 25:19]
  wire  d__GEN_437; // @[core.scala 25:19]
  wire  d__GEN_332_0; // @[core.scala 25:19]
  wire  d__GEN_126_1; // @[core.scala 25:19]
  wire  d__GEN_245_0; // @[core.scala 25:19]
  wire  d__GEN_359_0; // @[core.scala 25:19]
  wire  d__GEN_431; // @[core.scala 25:19]
  wire  d__GEN_458; // @[core.scala 25:19]
  wire  d__GEN_317_0; // @[core.scala 25:19]
  wire  d__GEN_326_0; // @[core.scala 25:19]
  wire  d__GEN_341_0; // @[core.scala 25:19]
  wire  d__GEN_1_3; // @[core.scala 25:19]
  wire  d__GEN_394_0; // @[core.scala 25:19]
  wire  d__GEN_248_0; // @[core.scala 25:19]
  wire  d__GEN_347_0; // @[core.scala 25:19]
  wire  d__GEN_92_1; // @[core.scala 25:19]
  wire  d__GEN_102_1; // @[core.scala 25:19]
  wire  d__GEN_425_0; // @[core.scala 25:19]
  wire  d__GEN_305_0; // @[core.scala 25:19]
  wire  d__GEN_419_0; // @[core.scala 25:19]
  wire  d__GEN_320_0; // @[core.scala 25:19]
  wire  d__GEN_108_1; // @[core.scala 25:19]
  wire  d__GEN_114_1; // @[core.scala 25:19]
  wire  d__GEN_123_1; // @[core.scala 25:19]
  wire  d__GEN_413_0; // @[core.scala 25:19]
  wire  d__GEN_440; // @[core.scala 25:19]
  wire  d__GEN_295_0; // @[core.scala 25:19]
  wire  d__GEN_129_1; // @[core.scala 25:19]
  wire  d__GEN_404_0; // @[core.scala 25:19]
  wire  d__GEN_403_0; // @[core.scala 25:19]
  wire  d__GEN_242_0; // @[core.scala 25:19]
  wire  d__GEN_15_1; // @[core.scala 25:19]
  wire  d__GEN_96_1; // @[core.scala 25:19]
  wire  d__GEN_86_1; // @[core.scala 25:19]
  wire  d__GEN_164_1; // @[core.scala 25:19]
  wire  d__GEN_308_0; // @[core.scala 25:19]
  wire  d__GEN_149_1; // @[core.scala 25:19]
  wire  d__GEN_329_0; // @[core.scala 25:19]
  wire  d__GEN_292_0; // @[core.scala 25:19]
  wire  d__GEN_298_0; // @[core.scala 25:19]
  wire  d__GEN_391_0; // @[core.scala 25:19]
  wire  d__GEN_314_0; // @[core.scala 25:19]
  wire  d__GEN_323_0; // @[core.scala 25:19]
  wire  d__GEN_376_0; // @[core.scala 25:19]
  wire  d__GEN_422_0; // @[core.scala 25:19]
  wire  d__GEN_277_0; // @[core.scala 25:19]
  wire  d__GEN_46_1; // @[core.scala 25:19]
  wire  d__GEN_111_1; // @[core.scala 25:19]
  wire  d__GEN_78_1; // @[core.scala 25:19]
  wire  d__GEN_407_0; // @[core.scala 25:19]
  wire  d__GEN_179_1; // @[core.scala 25:19]
  wire  d__GEN_397_0; // @[core.scala 25:19]
  wire  d__GEN_173_1; // @[core.scala 25:19]
  wire  d__GEN_70_1; // @[core.scala 25:19]
  wire  d__GEN_379_0; // @[core.scala 25:19]
  wire  d__GEN_82_1; // @[core.scala 25:19]
  wire  d__GEN_373_0; // @[core.scala 25:19]
  wire  d__GEN_54_1; // @[core.scala 25:19]
  wire  d__GEN_364_0; // @[core.scala 25:19]
  wire  d__GEN_259_0; // @[core.scala 25:19]
  wire  d__GEN_167_1; // @[core.scala 25:19]
  wire  d__GEN_43_1; // @[core.scala 25:19]
  wire  d__GEN_161_1; // @[core.scala 25:19]
  wire  d__GEN_265_0; // @[core.scala 25:19]
  wire  d__GEN_301_0; // @[core.scala 25:19]
  wire  d__GEN_146_2; // @[core.scala 25:19]
  wire  d__GEN_286_0; // @[core.scala 25:19]
  wire  d__GEN_400_0; // @[core.scala 25:19]
  wire  d__GEN_89_0; // @[core.scala 25:19]
  wire  d__GEN_358_0; // @[core.scala 25:19]
  wire  d__GEN_385_0; // @[core.scala 25:19]
  wire  d__GEN_457; // @[core.scala 25:19]
  wire  d__GEN_311_0; // @[core.scala 25:19]
  wire  d__GEN_280_0; // @[core.scala 25:19]
  wire  d__GEN_143_1; // @[core.scala 25:19]
  wire  d__GEN_367_0; // @[core.scala 25:19]
  wire  d__GEN_247_0; // @[core.scala 25:19]
  wire  d__GEN_274_0; // @[core.scala 25:19]
  wire  d__GEN_460; // @[core.scala 25:19]
  wire  d__GEN_283_0; // @[core.scala 25:19]
  wire  d__GEN_388_0; // @[core.scala 25:19]
  wire  d__GEN_382_0; // @[core.scala 25:19]
  wire  d__GEN_268_0; // @[core.scala 25:19]
  wire  d__GEN_176_1; // @[core.scala 25:19]
  wire  d__GEN_346_0; // @[core.scala 25:19]
  wire  d__GEN_64_1; // @[core.scala 25:19]
  wire  d__GEN_340_0; // @[core.scala 25:19]
  wire  d__GEN_134_1; // @[core.scala 25:19]
  wire  d__GEN_149_2; // @[core.scala 25:19]
  wire  d__GEN_439; // @[core.scala 25:19]
  wire  d__GEN_262_0; // @[core.scala 25:19]
  wire  d__GEN_17_1; // @[core.scala 25:19]
  wire  d__GEN_361_0; // @[core.scala 25:19]
  wire  d__GEN_155_1; // @[core.scala 25:19]
  wire  d__GEN_170_1; // @[core.scala 25:19]
  wire  d__GEN_73_1; // @[core.scala 25:19]
  wire  d__GEN_128_1; // @[core.scala 25:19]
  wire  d__GEN_241_0; // @[core.scala 25:19]
  wire  d__GEN_445; // @[core.scala 25:19]
  wire  d__GEN_289_0; // @[core.scala 25:19]
  wire  d__GEN_131_1; // @[core.scala 25:19]
  wire  d__GEN_152_2; // @[core.scala 25:19]
  wire  d__GEN_421_0; // @[core.scala 25:19]
  wire  d__GEN_427; // @[core.scala 25:19]
  wire  d__GEN_454; // @[core.scala 25:19]
  wire  d__GEN_256_0; // @[core.scala 25:19]
  wire  d__GEN_110_1; // @[core.scala 25:19]
  wire  d__GEN_40_1; // @[core.scala 25:19]
  wire  d__GEN_5_2; // @[core.scala 25:19]
  wire  d__GEN_158_1; // @[core.scala 25:19]
  wire  d__GEN_271_0; // @[core.scala 25:19]
  wire  d__GEN_322_0; // @[core.scala 25:19]
  wire  d__GEN_334_0; // @[core.scala 25:19]
  wire  d__GEN_116_1; // @[core.scala 25:19]
  wire  d__GEN_235_0; // @[core.scala 25:19]
  wire  d__GEN_349_0; // @[core.scala 25:19]
  wire  d__GEN_147_2; // @[core.scala 25:19]
  wire  d__GEN_448; // @[core.scala 25:19]
  wire  d__GEN_442; // @[core.scala 25:19]
  wire  d__GEN_343_0; // @[core.scala 25:19]
  wire  d__GEN_355_0; // @[core.scala 25:19]
  wire  d__GEN_137_1; // @[core.scala 25:19]
  wire  d__GEN_370_0; // @[core.scala 25:19]
  wire  d__GEN_250_0; // @[core.scala 25:19]
  wire  d__GEN_463; // @[core.scala 25:19]
  wire  d__GEN_328_0; // @[core.scala 25:19]
  CtlPath c ( // @[core.scala 24:19]
    .metaReset(c_metaReset),
    .clock(c_clock),
    .reset(c_reset),
    .io_imem_resp_valid(c_io_imem_resp_valid),
    .io_dmem_resp_valid(c_io_dmem_resp_valid),
    .io_dat_dec_inst(c_io_dat_dec_inst),
    .io_dat_exe_br_eq(c_io_dat_exe_br_eq),
    .io_dat_exe_br_lt(c_io_dat_exe_br_lt),
    .io_dat_exe_br_ltu(c_io_dat_exe_br_ltu),
    .io_dat_exe_br_type(c_io_dat_exe_br_type),
    .io_dat_mem_ctrl_dmem_val(c_io_dat_mem_ctrl_dmem_val),
    .io_dat_csr_eret(c_io_dat_csr_eret),
    .io_ctl_dec_stall(c_io_ctl_dec_stall),
    .io_ctl_full_stall(c_io_ctl_full_stall),
    .io_ctl_exe_pc_sel(c_io_ctl_exe_pc_sel),
    .io_ctl_br_type(c_io_ctl_br_type),
    .io_ctl_if_kill(c_io_ctl_if_kill),
    .io_ctl_dec_kill(c_io_ctl_dec_kill),
    .io_ctl_op1_sel(c_io_ctl_op1_sel),
    .io_ctl_op2_sel(c_io_ctl_op2_sel),
    .io_ctl_alu_fun(c_io_ctl_alu_fun),
    .io_ctl_wb_sel(c_io_ctl_wb_sel),
    .io_ctl_rf_wen(c_io_ctl_rf_wen),
    .io_ctl_mem_val(c_io_ctl_mem_val),
    .io_ctl_mem_fcn(c_io_ctl_mem_fcn),
    .io_ctl_mem_typ(c_io_ctl_mem_typ),
    .io_ctl_csr_cmd(c_io_ctl_csr_cmd),
    .io_ctl_fencei(c_io_ctl_fencei),
    .io_ctl_pipeline_kill(c_io_ctl_pipeline_kill),
    .io_ctl_mem_exception(c_io_ctl_mem_exception),
    ._GEN_111_0(c__GEN_111_0),
    ._GEN_71_0(c__GEN_71_0),
    ._GEN_324_0(c__GEN_324_0),
    ._GEN_219_0(c__GEN_219_0),
    ._GEN_168_0(c__GEN_168_0),
    ._GEN_1_0(c__GEN_1_0),
    ._GEN_423_0(c__GEN_423_0),
    ._GEN_44_0(c__GEN_44_0),
    ._GEN_267_0(c__GEN_267_0),
    ._GEN_126_0(c__GEN_126_0),
    ._GEN_153_0(c__GEN_153_0),
    ._GEN_225_0(c__GEN_225_0),
    ._GEN_59_0(c__GEN_59_0),
    ._GEN_252_0(c__GEN_252_0),
    ._GEN_147_0(c__GEN_147_0),
    ._GEN_351_0(c__GEN_351_0),
    ._GEN_210_0(c__GEN_210_0),
    ._GEN_246_0(c__GEN_246_0),
    ._GEN_65_0(c__GEN_65_0),
    ._GEN_132_0(c__GEN_132_0),
    ._GEN_318_0(c__GEN_318_0),
    ._GEN_92_0(c__GEN_92_0),
    ._GEN_345_0(c__GEN_345_0),
    ._GEN_231_0(c__GEN_231_0),
    ._GEN_417_0(c__GEN_417_0),
    ._GEN_50_0(c__GEN_50_0),
    ._GEN_330_0(c__GEN_330_0),
    ._GEN_86_0(c__GEN_86_0),
    ._GEN_339_0(c__GEN_339_0),
    ._GEN_240_0(c__GEN_240_0),
    ._GEN_234_0(c__GEN_234_0),
    ._GEN_120_0(c__GEN_120_0),
    ._GEN_129_0(c__GEN_129_0),
    ._GEN_333_0(c__GEN_333_0),
    ._GEN_302_0(c__GEN_302_0),
    ._GEN_228_0(c__GEN_228_0),
    ._GEN_197_0(c__GEN_197_0),
    ._GEN_411_0(c__GEN_411_0),
    ._GEN_401_0(c__GEN_401_0),
    ._GEN_47_0(c__GEN_47_0),
    ._GEN_296_0(c__GEN_296_0),
    ._GEN_74_0(c__GEN_74_0),
    ._GEN_213_0(c__GEN_213_0),
    ._GEN_32_0(c__GEN_32_0),
    ._GEN_68_0(c__GEN_68_0),
    ._GEN_135_0(c__GEN_135_0),
    ._GEN_26_0(c__GEN_26_0),
    ._GEN_53_0(c__GEN_53_0),
    ._GEN_141_0(c__GEN_141_0),
    ._GEN_327_0(c__GEN_327_0),
    ._GEN_395_0(c__GEN_395_0),
    ._GEN_249_0(c__GEN_249_0),
    ._GEN_114_0(c__GEN_114_0),
    ._GEN_312_0(c__GEN_312_0),
    ._GEN_203_0(c__GEN_203_0),
    ._GEN_20_0(c__GEN_20_0),
    ._GEN_15_0(c__GEN_15_0),
    ._GEN_216_0(c__GEN_216_0),
    ._GEN_206_0(c__GEN_206_0),
    ._GEN_420_0(c__GEN_420_0),
    ._GEN_123_0(c__GEN_123_0),
    ._GEN_315_0(c__GEN_315_0),
    ._GEN_284_0(c__GEN_284_0),
    ._GEN_179_0(c__GEN_179_0),
    ._GEN_222_0(c__GEN_222_0),
    ._GEN_377_0(c__GEN_377_0),
    ._GEN_191_0(c__GEN_191_0),
    ._GEN_290_0(c__GEN_290_0),
    ._GEN_404_0(c__GEN_404_0),
    ._GEN_56_1(c__GEN_56_1),
    ._GEN_305_0(c__GEN_305_0),
    ._GEN_299_0(c__GEN_299_0),
    ._GEN_185_0(c__GEN_185_0),
    ._GEN_398_0(c__GEN_398_0),
    ._GEN_41_0(c__GEN_41_0),
    ._GEN_321_0(c__GEN_321_0),
    ._GEN_414_0(c__GEN_414_0),
    ._GEN_383_0(c__GEN_383_0),
    ._GEN_35_0(c__GEN_35_0),
    ._GEN_29_0(c__GEN_29_0),
    ._GEN_278_0(c__GEN_278_0),
    ._GEN_117_0(c__GEN_117_0),
    ._GEN_365_0(c__GEN_365_0),
    ._GEN_359_0(c__GEN_359_0),
    ._GEN_38_0(c__GEN_38_0),
    ._GEN_167_0(c__GEN_167_0),
    ._GEN_350_0(c__GEN_350_0),
    ._GEN_106_0(c__GEN_106_0),
    ._GEN_18_0(c__GEN_18_0),
    ._GEN_293_0(c__GEN_293_0),
    ._GEN_371_0(c__GEN_371_0),
    ._GEN_251_0(c__GEN_251_0),
    ._GEN_209_0(c__GEN_209_0),
    ._GEN_308_0(c__GEN_308_0),
    ._GEN_173_0(c__GEN_173_0),
    ._GEN_200_0(c__GEN_200_0),
    ._GEN_386_0(c__GEN_386_0),
    ._GEN_272_0(c__GEN_272_0),
    ._GEN_91_1(c__GEN_91_1),
    ._GEN_194_0(c__GEN_194_0),
    ._GEN_188_0(c__GEN_188_0),
    ._GEN_392_0(c__GEN_392_0),
    ._GEN_23_0(c__GEN_23_0),
    ._GEN_407_0(c__GEN_407_0),
    ._GEN_287_0(c__GEN_287_0),
    ._GEN_266_0(c__GEN_266_0),
    ._GEN_374_0(c__GEN_374_0),
    ._GEN_233_0(c__GEN_233_0),
    ._GEN_269_0(c__GEN_269_0),
    ._GEN_260_0(c__GEN_260_0),
    ._GEN_161_0(c__GEN_161_0),
    ._GEN_155_0(c__GEN_155_0),
    ._GEN_368_0(c__GEN_368_0),
    ._GEN_254_0(c__GEN_254_0),
    ._GEN_281_0(c__GEN_281_0),
    ._GEN_73_0(c__GEN_73_0),
    ._GEN_353_0(c__GEN_353_0),
    ._GEN_332_0(c__GEN_332_0),
    ._GEN_88_1(c__GEN_88_1),
    ._GEN_176_0(c__GEN_176_0),
    ._GEN_380_0(c__GEN_380_0),
    ._GEN_389_0(c__GEN_389_0),
    ._GEN_94_0(c__GEN_94_0),
    ._GEN_347_0(c__GEN_347_0),
    ._GEN_109_0(c__GEN_109_0),
    ._GEN_182_0(c__GEN_182_0),
    ._GEN_9_0(c__GEN_9_0),
    ._GEN_149_0(c__GEN_149_0),
    ._GEN_248_0(c__GEN_248_0),
    ._GEN_275_0(c__GEN_275_0),
    ._GEN_140_1(c__GEN_140_1),
    ._GEN_100_0(c__GEN_100_0),
    ._GEN_362_0(c__GEN_362_0),
    ._GEN_413_0(c__GEN_413_0),
    ._GEN_76_0(c__GEN_76_0),
    ._GEN_164_0(c__GEN_164_0),
    ._GEN_242_0(c__GEN_242_0),
    ._GEN_137_0(c__GEN_137_0),
    ._GEN_341_0(c__GEN_341_0),
    ._GEN_263_0(c__GEN_263_0),
    ._GEN_257_0(c__GEN_257_0),
    ._GEN_122_1(c__GEN_122_1),
    ._GEN_143_0(c__GEN_143_0),
    ._GEN_82_0(c__GEN_82_0),
    ._GEN_170_0(c__GEN_170_0),
    ._GEN_356_0(c__GEN_356_0),
    ._GEN_221_0(c__GEN_221_0),
    ._GEN_215_0(c__GEN_215_0),
    ._GEN_320_0(c__GEN_320_0),
    ._GEN_314_0(c__GEN_314_0),
    ._GEN_329_0(c__GEN_329_0),
    ._GEN_103_1(c__GEN_103_1),
    ._GEN_97_0(c__GEN_97_0),
    ._GEN_236_0(c__GEN_236_0),
    ._GEN_61_0(c__GEN_61_0),
    ._GEN_55_0(c__GEN_55_0),
    ._GEN_335_0(c__GEN_335_0),
    ._GEN_158_0(c__GEN_158_0),
    ._GEN_422_0(c__GEN_422_0),
    ._GEN_245_0(c__GEN_245_0),
    ._GEN_37_0(c__GEN_37_0),
    ._GEN_125_1(c__GEN_125_1),
    ._GEN_70_0(c__GEN_70_0),
    ._GEN_64_0(c__GEN_64_0),
    ._GEN_344_0(c__GEN_344_0),
    ._GEN_338_0(c__GEN_338_0),
    ._GEN_416_0(c__GEN_416_0),
    ._GEN_406_1(c__GEN_406_1),
    ._GEN_58_0(c__GEN_58_0),
    ._GEN_85_1(c__GEN_85_1),
    ._GEN_43_0(c__GEN_43_0),
    ._GEN_131_0(c__GEN_131_0),
    ._GEN_230_0(c__GEN_230_0),
    ._GEN_239_0(c__GEN_239_0),
    ._GEN_152_0(c__GEN_152_0),
    ._GEN_307_1(c__GEN_307_1),
    ._GEN_146_1(c__GEN_146_1),
    ._GEN_224_0(c__GEN_224_0),
    ._GEN_110_0(c__GEN_110_0),
    ._GEN_119_1(c__GEN_119_1),
    ._GEN_323_0(c__GEN_323_0),
    ._GEN_317_0(c__GEN_317_0),
    ._GEN_79_1(c__GEN_79_1),
    ._GEN_218_0(c__GEN_218_0),
    ._GEN_208_0(c__GEN_208_0),
    ._GEN_196_0(c__GEN_196_0),
    ._GEN_31_0(c__GEN_31_0),
    ._GEN_400_0(c__GEN_400_0),
    ._GEN_113_1(c__GEN_113_1),
    ._GEN_212_0(c__GEN_212_0),
    ._GEN_181_0(c__GEN_181_0),
    ._GEN_227_0(c__GEN_227_0),
    ._GEN_425_0(c__GEN_425_0),
    ._GEN_280_0(c__GEN_280_0),
    ._GEN_46_0(c__GEN_46_0),
    ._GEN_134_0(c__GEN_134_0),
    ._GEN_289_0(c__GEN_289_0),
    ._GEN_202_0(c__GEN_202_0),
    ._GEN_419_0(c__GEN_419_0),
    ._GEN_388_0(c__GEN_388_0),
    ._GEN_410_0(c__GEN_410_0),
    ._GEN_52_0(c__GEN_52_0),
    ._GEN_311_0(c__GEN_311_0),
    ._GEN_301_0(c__GEN_301_0),
    ._GEN_295_0(c__GEN_295_0),
    ._GEN_67_0(c__GEN_67_0),
    ._GEN_25_0(c__GEN_25_0),
    ._GEN_409_1(c__GEN_409_1),
    ._GEN_326_0(c__GEN_326_0),
    ._GEN_394_0(c__GEN_394_0),
    ._GEN_128_0(c__GEN_128_0),
    ._GEN_376_0(c__GEN_376_0),
    ._GEN_40_0(c__GEN_40_0),
    ._GEN_34_0(c__GEN_34_0),
    ._GEN_49_0(c__GEN_49_0),
    ._GEN_102_0(c__GEN_102_0),
    ._GEN_190_0(c__GEN_190_0),
    ._GEN_205_0(c__GEN_205_0),
    ._GEN_298_0(c__GEN_298_0),
    ._GEN_163_1(c__GEN_163_1),
    ._GEN_14_0(c__GEN_14_0),
    ._GEN_116_0(c__GEN_116_0),
    ._GEN_283_0(c__GEN_283_0),
    ._GEN_184_0(c__GEN_184_0),
    ._GEN_178_1(c__GEN_178_1),
    ._GEN_382_0(c__GEN_382_0),
    ._GEN_397_0(c__GEN_397_0),
    ._GEN_277_0(c__GEN_277_0),
    ._GEN_304_1(c__GEN_304_1),
    ._GEN_199_0(c__GEN_199_0),
    ._GEN_403_0(c__GEN_403_0),
    ._GEN_262_0(c__GEN_262_0),
    ._GEN_28_0(c__GEN_28_0),
    ._GEN_361_0(c__GEN_361_0),
    ._GEN_96_0(c__GEN_96_0),
    ._GEN_193_0(c__GEN_193_0),
    ._GEN_379_0(c__GEN_379_0),
    ._GEN_244_1(c__GEN_244_1),
    ._GEN_271_0(c__GEN_271_0),
    ._GEN_151_2(c__GEN_151_2),
    ._GEN_166_1(c__GEN_166_1),
    ._GEN_370_0(c__GEN_370_0),
    ._GEN_364_0(c__GEN_364_0),
    ._GEN_259_0(c__GEN_259_0),
    ._GEN_292_0(c__GEN_292_0),
    ._GEN_84_0(c__GEN_84_0),
    ._GEN_78_0(c__GEN_78_0),
    ._GEN_385_0(c__GEN_385_0),
    ._GEN_250_0(c__GEN_250_0),
    ._GEN_343_0(c__GEN_343_0),
    ._GEN_105_0(c__GEN_105_0),
    ._GEN_99_0(c__GEN_99_0),
    ._GEN_358_0(c__GEN_358_0),
    ._GEN_22_0(c__GEN_22_0),
    ._GEN_265_0(c__GEN_265_0),
    ._GEN_17_0(c__GEN_17_0),
    ._GEN_90_1(c__GEN_90_1),
    ._GEN_172_1(c__GEN_172_1),
    ._GEN_187_0(c__GEN_187_0),
    ._GEN_391_0(c__GEN_391_0),
    ._GEN_286_0(c__GEN_286_0),
    ._GEN_145_1(c__GEN_145_1),
    ._GEN_232_0(c__GEN_232_0),
    ._GEN_274_0(c__GEN_274_0),
    ._GEN_175_1(c__GEN_175_1),
    ._GEN_169_1(c__GEN_169_1),
    ._GEN_247_0(c__GEN_247_0),
    ._GEN_133_1(c__GEN_133_1),
    ._GEN_160_1(c__GEN_160_1),
    ._GEN_346_0(c__GEN_346_0),
    ._GEN_373_0(c__GEN_373_0),
    ._GEN_424_1(c__GEN_424_1),
    ._GEN_268_0(c__GEN_268_0),
    ._GEN_127_1(c__GEN_127_1),
    ._GEN_8_0(c__GEN_8_0),
    ._GEN_331_1(c__GEN_331_1),
    ._GEN_93_1(c__GEN_93_1),
    ._GEN_87_1(c__GEN_87_1),
    ._GEN_367_0(c__GEN_367_0),
    ._GEN_226_0(c__GEN_226_0),
    ._GEN_253_1(c__GEN_253_1),
    ._GEN_325_1(c__GEN_325_1),
    ._GEN_148_1(c__GEN_148_1),
    ._GEN_352_1(c__GEN_352_1),
    ._GEN_108_0(c__GEN_108_0),
    ._GEN_72_1(c__GEN_72_1),
    ._GEN_66_0(c__GEN_66_0),
    ._GEN_154_1(c__GEN_154_1),
    ._GEN_241_0(c__GEN_241_0),
    ._GEN_402_1(c__GEN_402_1),
    ._GEN_48_0(c__GEN_48_0),
    ._GEN_60_0(c__GEN_60_0),
    ._GEN_75_1(c__GEN_75_1),
    ._GEN_349_0(c__GEN_349_0),
    ._GEN_214_0(c__GEN_214_0),
    ._GEN_412_1(c__GEN_412_1),
    ._GEN_256_0(c__GEN_256_0),
    ._GEN_121_1(c__GEN_121_1),
    ._GEN_81_0(c__GEN_81_0),
    ._GEN_54_0(c__GEN_54_0),
    ._GEN_136_1(c__GEN_136_1),
    ._GEN_142_1(c__GEN_142_1),
    ._GEN_340_0(c__GEN_340_0),
    ._GEN_355_0(c__GEN_355_0),
    ._GEN_235_0(c__GEN_235_0),
    ._GEN_313_1(c__GEN_313_1),
    ._GEN_69_1(c__GEN_69_1),
    ._GEN_157_1(c__GEN_157_1),
    ._GEN_220_0(c__GEN_220_0),
    ._GEN_229_0(c__GEN_229_0),
    ._GEN_115_1(c__GEN_115_1),
    ._GEN_334_0(c__GEN_334_0),
    ._GEN_328_0(c__GEN_328_0),
    ._GEN_36_0(c__GEN_36_0),
    ._GEN_405_1(c__GEN_405_1),
    ._GEN_415_1(c__GEN_415_1),
    ._GEN_124_1(c__GEN_124_1),
    ._GEN_322_0(c__GEN_322_0),
    ._GEN_337_1(c__GEN_337_1),
    ._GEN_223_0(c__GEN_223_0),
    ._GEN_217_0(c__GEN_217_0),
    ._GEN_192_0(c__GEN_192_0),
    ._GEN_390_1(c__GEN_390_1),
    ._GEN_42_1(c__GEN_42_1),
    ._GEN_291_1(c__GEN_291_1),
    ._GEN_139_1(c__GEN_139_1),
    ._GEN_207_0(c__GEN_207_0),
    ._GEN_399_1(c__GEN_399_1),
    ._GEN_421_0(c__GEN_421_0),
    ._GEN_63_0(c__GEN_63_0),
    ._GEN_316_1(c__GEN_316_1),
    ._GEN_306_1(c__GEN_306_1),
    ._GEN_21_1(c__GEN_21_1),
    ._GEN_384_1(c__GEN_384_1),
    ._GEN_118_1(c__GEN_118_1),
    ._GEN_57_0(c__GEN_57_0),
    ._GEN_130_1(c__GEN_130_1),
    ._GEN_238_1(c__GEN_238_1),
    ._GEN_45_1(c__GEN_45_1),
    ._GEN_201_0(c__GEN_201_0),
    ._GEN_195_0(c__GEN_195_0),
    ._GEN_309_1(c__GEN_309_1),
    ._GEN_372_1(c__GEN_372_1),
    ._GEN_19_0(c__GEN_19_0),
    ._GEN_51_0(c__GEN_51_0),
    ._GEN_294_1(c__GEN_294_1),
    ._GEN_180_0(c__GEN_180_0),
    ._GEN_189_0(c__GEN_189_0),
    ._GEN_211_0(c__GEN_211_0),
    ._GEN_393_1(c__GEN_393_1),
    ._GEN_387_1(c__GEN_387_1),
    ._GEN_39_0(c__GEN_39_0),
    ._GEN_288_1(c__GEN_288_1),
    ._GEN_310_1(c__GEN_310_1),
    ._GEN_300_1(c__GEN_300_1),
    ._GEN_319_1(c__GEN_319_1),
    ._GEN_107_1(c__GEN_107_1),
    ._GEN_174_1(c__GEN_174_1),
    ._GEN_30_0(c__GEN_30_0),
    ._GEN_24_0(c__GEN_24_0),
    ._GEN_408_1(c__GEN_408_1),
    ._GEN_418_1(c__GEN_418_1),
    ._GEN_273_1(c__GEN_273_1),
    ._GEN_5_1(c__GEN_5_1),
    ._GEN_112_1(c__GEN_112_1),
    ._GEN_366_1(c__GEN_366_1),
    ._GEN_360_1(c__GEN_360_1),
    ._GEN_354_1(c__GEN_354_1),
    ._GEN_33_1(c__GEN_33_1),
    ._GEN_276_1(c__GEN_276_1),
    ._GEN_348_1(c__GEN_348_1),
    ._GEN_101_1(c__GEN_101_1),
    ._GEN_375_1(c__GEN_375_1),
    ._GEN_27_0(c__GEN_27_0),
    ._GEN_13_0(c__GEN_13_0),
    ._GEN_297_1(c__GEN_297_1),
    ._GEN_89_1(c__GEN_89_1),
    ._GEN_177_1(c__GEN_177_1),
    ._GEN_255_1(c__GEN_255_1),
    ._GEN_204_0(c__GEN_204_0),
    ._GEN_80_1(c__GEN_80_1),
    ._GEN_303_1(c__GEN_303_1),
    ._GEN_162_1(c__GEN_162_1),
    ._GEN_198_0(c__GEN_198_0),
    ._GEN_381_1(c__GEN_381_1),
    ._GEN_261_1(c__GEN_261_1),
    ._GEN_156_1(c__GEN_156_1),
    ._GEN_95_1(c__GEN_95_1),
    ._GEN_183_0(c__GEN_183_0),
    ._GEN_369_1(c__GEN_369_1),
    ._GEN_282_1(c__GEN_282_1),
    ._GEN_396_1(c__GEN_396_1),
    ._GEN_378_1(c__GEN_378_1),
    ._GEN_186_0(c__GEN_186_0),
    ._GEN_62_0(c__GEN_62_0),
    ._GEN_285_1(c__GEN_285_1),
    ._GEN_336_1(c__GEN_336_1),
    ._GEN_144_1(c__GEN_144_1),
    ._GEN_150_2(c__GEN_150_2),
    ._GEN_363_1(c__GEN_363_1),
    ._GEN_243_1(c__GEN_243_1),
    ._GEN_258_1(c__GEN_258_1),
    ._GEN_138_1(c__GEN_138_1),
    ._GEN_171_1(c__GEN_171_1),
    ._GEN_357_1(c__GEN_357_1),
    ._GEN_165_1(c__GEN_165_1),
    ._GEN_264_1(c__GEN_264_1),
    ._GEN_16_1(c__GEN_16_1),
    ._GEN_342_1(c__GEN_342_1),
    ._GEN_98_1(c__GEN_98_1),
    ._GEN_237_1(c__GEN_237_1),
    ._GEN_83_1(c__GEN_83_1),
    ._GEN_77_0(c__GEN_77_0),
    ._GEN_270_1(c__GEN_270_1),
    ._GEN_279_1(c__GEN_279_1),
    ._GEN_159_1(c__GEN_159_1),
    ._GEN_104_1(c__GEN_104_1)
  );
  DatPath d ( // @[core.scala 25:19]
    .metaReset(d_metaReset),
    .clock(d_clock),
    .reset(d_reset),
    .io_imem_req_bits_addr(d_io_imem_req_bits_addr),
    .io_imem_resp_bits_data(d_io_imem_resp_bits_data),
    .io_dmem_req_valid(d_io_dmem_req_valid),
    .io_dmem_req_bits_addr(d_io_dmem_req_bits_addr),
    .io_dmem_req_bits_data(d_io_dmem_req_bits_data),
    .io_dmem_req_bits_fcn(d_io_dmem_req_bits_fcn),
    .io_dmem_req_bits_typ(d_io_dmem_req_bits_typ),
    .io_dmem_resp_bits_data(d_io_dmem_resp_bits_data),
    .io_ctl_dec_stall(d_io_ctl_dec_stall),
    .io_ctl_full_stall(d_io_ctl_full_stall),
    .io_ctl_exe_pc_sel(d_io_ctl_exe_pc_sel),
    .io_ctl_br_type(d_io_ctl_br_type),
    .io_ctl_if_kill(d_io_ctl_if_kill),
    .io_ctl_dec_kill(d_io_ctl_dec_kill),
    .io_ctl_op1_sel(d_io_ctl_op1_sel),
    .io_ctl_op2_sel(d_io_ctl_op2_sel),
    .io_ctl_alu_fun(d_io_ctl_alu_fun),
    .io_ctl_wb_sel(d_io_ctl_wb_sel),
    .io_ctl_rf_wen(d_io_ctl_rf_wen),
    .io_ctl_mem_val(d_io_ctl_mem_val),
    .io_ctl_mem_fcn(d_io_ctl_mem_fcn),
    .io_ctl_mem_typ(d_io_ctl_mem_typ),
    .io_ctl_csr_cmd(d_io_ctl_csr_cmd),
    .io_ctl_fencei(d_io_ctl_fencei),
    .io_ctl_pipeline_kill(d_io_ctl_pipeline_kill),
    .io_ctl_mem_exception(d_io_ctl_mem_exception),
    .io_dat_dec_inst(d_io_dat_dec_inst),
    .io_dat_exe_br_eq(d_io_dat_exe_br_eq),
    .io_dat_exe_br_lt(d_io_dat_exe_br_lt),
    .io_dat_exe_br_ltu(d_io_dat_exe_br_ltu),
    .io_dat_exe_br_type(d_io_dat_exe_br_type),
    .io_dat_mem_ctrl_dmem_val(d_io_dat_mem_ctrl_dmem_val),
    .io_dat_csr_eret(d_io_dat_csr_eret),
    ._GEN_451(d__GEN_451),
    ._GEN_331(d__GEN_331),
    ._GEN_337(d__GEN_337),
    ._GEN_113_0(d__GEN_113_0),
    ._GEN_415(d__GEN_415),
    ._GEN_436(d__GEN_436),
    ._GEN_140_0(d__GEN_140_0),
    ._GEN_98_0(d__GEN_98_0),
    ._GEN_352(d__GEN_352),
    ._GEN_125_0(d__GEN_125_0),
    ._GEN_430(d__GEN_430),
    ._GEN_119_0(d__GEN_119_0),
    ._GEN_88_0(d__GEN_88_0),
    ._GEN_151_0(d__GEN_151_0),
    ._GEN_310(d__GEN_310),
    ._GEN_104_0(d__GEN_104_0),
    ._GEN_409(d__GEN_409),
    ._GEN_253(d__GEN_253),
    ._GEN_316(d__GEN_316),
    ._GEN_244(d__GEN_244),
    ._GEN_238(d__GEN_238),
    ._GEN_101_0(d__GEN_101_0),
    ._GEN_325(d__GEN_325),
    ._GEN_169_0(d__GEN_169_0),
    ._GEN_433(d__GEN_433),
    ._GEN_313(d__GEN_313),
    ._GEN_91_0(d__GEN_91_0),
    ._GEN_11_0(d__GEN_11_0),
    ._GEN_304(d__GEN_304),
    ._GEN_294(d__GEN_294),
    ._GEN_303(d__GEN_303),
    ._GEN_107_0(d__GEN_107_0),
    ._GEN_0_0(d__GEN_0_0),
    ._GEN_402(d__GEN_402),
    ._GEN_412(d__GEN_412),
    ._GEN_424(d__GEN_424),
    ._GEN_175_0(d__GEN_175_0),
    ._GEN_319(d__GEN_319),
    ._GEN_288(d__GEN_288),
    ._GEN_56_0(d__GEN_56_0),
    ._GEN_418(d__GEN_418),
    ._GEN_122_0(d__GEN_122_0),
    ._GEN_387(d__GEN_387),
    ._GEN_72_0(d__GEN_72_0),
    ._GEN_75_0(d__GEN_75_0),
    ._GEN_85_0(d__GEN_85_0),
    ._GEN_178_0(d__GEN_178_0),
    ._GEN_157_0(d__GEN_157_0),
    ._GEN_462(d__GEN_462),
    ._GEN_69_0(d__GEN_69_0),
    ._GEN_375(d__GEN_375),
    ._GEN_151_1(d__GEN_151_1),
    ._GEN_33_0(d__GEN_33_0),
    ._GEN_390(d__GEN_390),
    ._GEN_307(d__GEN_307),
    ._GEN_297(d__GEN_297),
    ._GEN_406(d__GEN_406),
    ._GEN_270(d__GEN_270),
    ._GEN_95_0(d__GEN_95_0),
    ._GEN_45_0(d__GEN_45_0),
    ._GEN_369(d__GEN_369),
    ._GEN_396(d__GEN_396),
    ._GEN_172_0(d__GEN_172_0),
    ._GEN_276(d__GEN_276),
    ._GEN_291(d__GEN_291),
    ._GEN_258(d__GEN_258),
    ._GEN_372(d__GEN_372),
    ._GEN_252_0(d__GEN_252_0),
    ._GEN_166_0(d__GEN_166_0),
    ._GEN_285(d__GEN_285),
    ._GEN_42_0(d__GEN_42_0),
    ._GEN_384(d__GEN_384),
    ._GEN_378(d__GEN_378),
    ._GEN_393(d__GEN_393),
    ._GEN_273(d__GEN_273),
    ._GEN_456(d__GEN_456),
    ._GEN_80_0(d__GEN_80_0),
    ._GEN_351_0(d__GEN_351_0),
    ._GEN_139_0(d__GEN_139_0),
    ._GEN_145_0(d__GEN_145_0),
    ._GEN_450(d__GEN_450),
    ._GEN_53_1(d__GEN_53_1),
    ._GEN_357(d__GEN_357),
    ._GEN_160_0(d__GEN_160_0),
    ._GEN_279(d__GEN_279),
    ._GEN_133_0(d__GEN_133_0),
    ._GEN_399(d__GEN_399),
    ._GEN_264(d__GEN_264),
    ._GEN_300(d__GEN_300),
    ._GEN_127_0(d__GEN_127_0),
    ._GEN_432(d__GEN_432),
    ._GEN_381(d__GEN_381),
    ._GEN_339_0(d__GEN_339_0),
    ._GEN_261(d__GEN_261),
    ._GEN_16_0(d__GEN_16_0),
    ._GEN_360(d__GEN_360),
    ._GEN_163_0(d__GEN_163_0),
    ._GEN_246_0(d__GEN_246_0),
    ._GEN_438(d__GEN_438),
    ._GEN_282(d__GEN_282),
    ._GEN_345_0(d__GEN_345_0),
    ._GEN_121_0(d__GEN_121_0),
    ._GEN_240_0(d__GEN_240_0),
    ._GEN_148_0(d__GEN_148_0),
    ._GEN_154_0(d__GEN_154_0),
    ._GEN_444(d__GEN_444),
    ._GEN_267_0(d__GEN_267_0),
    ._GEN_459(d__GEN_459),
    ._GEN_453(d__GEN_453),
    ._GEN_366(d__GEN_366),
    ._GEN_7_0(d__GEN_7_0),
    ._GEN_142_0(d__GEN_142_0),
    ._GEN_324_0(d__GEN_324_0),
    ._GEN_333_0(d__GEN_333_0),
    ._GEN_342(d__GEN_342),
    ._GEN_405(d__GEN_405),
    ._GEN_420_0(d__GEN_420_0),
    ._GEN_306(d__GEN_306),
    ._GEN_109_1(d__GEN_109_1),
    ._GEN_103_0(d__GEN_103_0),
    ._GEN_3_0(d__GEN_3_0),
    ._GEN_136_0(d__GEN_136_0),
    ._GEN_426(d__GEN_426),
    ._GEN_441(d__GEN_441),
    ._GEN_94_1(d__GEN_94_1),
    ._GEN_348(d__GEN_348),
    ._GEN_255(d__GEN_255),
    ._GEN_115_0(d__GEN_115_0),
    ._GEN_146_0(d__GEN_146_0),
    ._GEN_363(d__GEN_363),
    ._GEN_321_0(d__GEN_321_0),
    ._GEN_327_0(d__GEN_327_0),
    ._GEN_354(d__GEN_354),
    ._GEN_234_0(d__GEN_234_0),
    ._GEN_130_0(d__GEN_130_0),
    ._GEN_249_0(d__GEN_249_0),
    ._GEN_243(d__GEN_243),
    ._GEN_447(d__GEN_447),
    ._GEN_330_0(d__GEN_330_0),
    ._GEN_429(d__GEN_429),
    ._GEN_293_0(d__GEN_293_0),
    ._GEN_87_0(d__GEN_87_0),
    ._GEN_414_0(d__GEN_414_0),
    ._GEN_309(d__GEN_309),
    ._GEN_299_0(d__GEN_299_0),
    ._GEN_336(d__GEN_336),
    ._GEN_408(d__GEN_408),
    ._GEN_112_0(d__GEN_112_0),
    ._GEN_150_0(d__GEN_150_0),
    ._GEN_435(d__GEN_435),
    ._GEN_97_1(d__GEN_97_1),
    ._GEN_124_0(d__GEN_124_0),
    ._GEN_118_0(d__GEN_118_0),
    ._GEN_392_0(d__GEN_392_0),
    ._GEN_398_0(d__GEN_398_0),
    ._GEN_423_0(d__GEN_423_0),
    ._GEN_237(d__GEN_237),
    ._GEN_315_0(d__GEN_315_0),
    ._GEN_79_0(d__GEN_79_0),
    ._GEN_1_2(d__GEN_1_2),
    ._GEN_90_0(d__GEN_90_0),
    ._GEN_162_0(d__GEN_162_0),
    ._GEN_302_0(d__GEN_302_0),
    ._GEN_106_1(d__GEN_106_1),
    ._GEN_71_1(d__GEN_71_1),
    ._GEN_380_0(d__GEN_380_0),
    ._GEN_174_0(d__GEN_174_0),
    ._GEN_318_0(d__GEN_318_0),
    ._GEN_287_0(d__GEN_287_0),
    ._GEN_386_0(d__GEN_386_0),
    ._GEN_281_0(d__GEN_281_0),
    ._GEN_312_0(d__GEN_312_0),
    ._GEN_417_0(d__GEN_417_0),
    ._GEN_411_0(d__GEN_411_0),
    ._GEN_55_1(d__GEN_55_1),
    ._GEN_100_1(d__GEN_100_1),
    ._GEN_168_1(d__GEN_168_1),
    ._GEN_401_0(d__GEN_401_0),
    ._GEN_44_1(d__GEN_44_1),
    ._GEN_74_1(d__GEN_74_1),
    ._GEN_374_0(d__GEN_374_0),
    ._GEN_368_0(d__GEN_368_0),
    ._GEN_383_0(d__GEN_383_0),
    ._GEN_263_0(d__GEN_263_0),
    ._GEN_177_0(d__GEN_177_0),
    ._GEN_171_0(d__GEN_171_0),
    ._GEN_446(d__GEN_446),
    ._GEN_290_0(d__GEN_290_0),
    ._GEN_83_0(d__GEN_83_0),
    ._GEN_135_1(d__GEN_135_1),
    ._GEN_389_0(d__GEN_389_0),
    ._GEN_93_0(d__GEN_93_0),
    ._GEN_254_0(d__GEN_254_0),
    ._GEN_21_0(d__GEN_21_0),
    ._GEN_461(d__GEN_461),
    ._GEN_362_0(d__GEN_362_0),
    ._GEN_156_0(d__GEN_156_0),
    ._GEN_150_1(d__GEN_150_1),
    ._GEN_68_1(d__GEN_68_1),
    ._GEN_296_0(d__GEN_296_0),
    ._GEN_395_0(d__GEN_395_0),
    ._GEN_275_0(d__GEN_275_0),
    ._GEN_269_0(d__GEN_269_0),
    ._GEN_278_0(d__GEN_278_0),
    ._GEN_138_0(d__GEN_138_0),
    ._GEN_251_0(d__GEN_251_0),
    ._GEN_455(d__GEN_455),
    ._GEN_377_0(d__GEN_377_0),
    ._GEN_153_1(d__GEN_153_1),
    ._GEN_272_0(d__GEN_272_0),
    ._GEN_47_1(d__GEN_47_1),
    ._GEN_335_0(d__GEN_335_0),
    ._GEN_41_1(d__GEN_41_1),
    ._GEN_434(d__GEN_434),
    ._GEN_257_0(d__GEN_257_0),
    ._GEN_443(d__GEN_443),
    ._GEN_356_0(d__GEN_356_0),
    ._GEN_350_0(d__GEN_350_0),
    ._GEN_132_1(d__GEN_132_1),
    ._GEN_144_0(d__GEN_144_0),
    ._GEN_159_0(d__GEN_159_0),
    ._GEN_428(d__GEN_428),
    ._GEN_449(d__GEN_449),
    ._GEN_117_1(d__GEN_117_1),
    ._GEN_236_0(d__GEN_236_0),
    ._GEN_371_0(d__GEN_371_0),
    ._GEN_165_0(d__GEN_165_0),
    ._GEN_284_0(d__GEN_284_0),
    ._GEN_147_1(d__GEN_147_1),
    ._GEN_416_0(d__GEN_416_0),
    ._GEN_260_0(d__GEN_260_0),
    ._GEN_105_1(d__GEN_105_1),
    ._GEN_338_0(d__GEN_338_0),
    ._GEN_141_1(d__GEN_141_1),
    ._GEN_99_1(d__GEN_99_1),
    ._GEN_344_0(d__GEN_344_0),
    ._GEN_239_0(d__GEN_239_0),
    ._GEN_353_0(d__GEN_353_0),
    ._GEN_266_0(d__GEN_266_0),
    ._GEN_452(d__GEN_452),
    ._GEN_120_1(d__GEN_120_1),
    ._GEN_365_0(d__GEN_365_0),
    ._GEN_6_0(d__GEN_6_0),
    ._GEN_410_0(d__GEN_410_0),
    ._GEN_152_1(d__GEN_152_1),
    ._GEN_437(d__GEN_437),
    ._GEN_332_0(d__GEN_332_0),
    ._GEN_126_1(d__GEN_126_1),
    ._GEN_245_0(d__GEN_245_0),
    ._GEN_359_0(d__GEN_359_0),
    ._GEN_431(d__GEN_431),
    ._GEN_458(d__GEN_458),
    ._GEN_317_0(d__GEN_317_0),
    ._GEN_326_0(d__GEN_326_0),
    ._GEN_341_0(d__GEN_341_0),
    ._GEN_1_3(d__GEN_1_3),
    ._GEN_394_0(d__GEN_394_0),
    ._GEN_248_0(d__GEN_248_0),
    ._GEN_347_0(d__GEN_347_0),
    ._GEN_92_1(d__GEN_92_1),
    ._GEN_102_1(d__GEN_102_1),
    ._GEN_425_0(d__GEN_425_0),
    ._GEN_305_0(d__GEN_305_0),
    ._GEN_419_0(d__GEN_419_0),
    ._GEN_320_0(d__GEN_320_0),
    ._GEN_108_1(d__GEN_108_1),
    ._GEN_114_1(d__GEN_114_1),
    ._GEN_123_1(d__GEN_123_1),
    ._GEN_413_0(d__GEN_413_0),
    ._GEN_440(d__GEN_440),
    ._GEN_295_0(d__GEN_295_0),
    ._GEN_129_1(d__GEN_129_1),
    ._GEN_404_0(d__GEN_404_0),
    ._GEN_403_0(d__GEN_403_0),
    ._GEN_242_0(d__GEN_242_0),
    ._GEN_15_1(d__GEN_15_1),
    ._GEN_96_1(d__GEN_96_1),
    ._GEN_86_1(d__GEN_86_1),
    ._GEN_164_1(d__GEN_164_1),
    ._GEN_308_0(d__GEN_308_0),
    ._GEN_149_1(d__GEN_149_1),
    ._GEN_329_0(d__GEN_329_0),
    ._GEN_292_0(d__GEN_292_0),
    ._GEN_298_0(d__GEN_298_0),
    ._GEN_391_0(d__GEN_391_0),
    ._GEN_314_0(d__GEN_314_0),
    ._GEN_323_0(d__GEN_323_0),
    ._GEN_376_0(d__GEN_376_0),
    ._GEN_422_0(d__GEN_422_0),
    ._GEN_277_0(d__GEN_277_0),
    ._GEN_46_1(d__GEN_46_1),
    ._GEN_111_1(d__GEN_111_1),
    ._GEN_78_1(d__GEN_78_1),
    ._GEN_407_0(d__GEN_407_0),
    ._GEN_179_1(d__GEN_179_1),
    ._GEN_397_0(d__GEN_397_0),
    ._GEN_173_1(d__GEN_173_1),
    ._GEN_70_1(d__GEN_70_1),
    ._GEN_379_0(d__GEN_379_0),
    ._GEN_82_1(d__GEN_82_1),
    ._GEN_373_0(d__GEN_373_0),
    ._GEN_54_1(d__GEN_54_1),
    ._GEN_364_0(d__GEN_364_0),
    ._GEN_259_0(d__GEN_259_0),
    ._GEN_167_1(d__GEN_167_1),
    ._GEN_43_1(d__GEN_43_1),
    ._GEN_161_1(d__GEN_161_1),
    ._GEN_265_0(d__GEN_265_0),
    ._GEN_301_0(d__GEN_301_0),
    ._GEN_146_2(d__GEN_146_2),
    ._GEN_286_0(d__GEN_286_0),
    ._GEN_400_0(d__GEN_400_0),
    ._GEN_89_0(d__GEN_89_0),
    ._GEN_358_0(d__GEN_358_0),
    ._GEN_385_0(d__GEN_385_0),
    ._GEN_457(d__GEN_457),
    ._GEN_311_0(d__GEN_311_0),
    ._GEN_280_0(d__GEN_280_0),
    ._GEN_143_1(d__GEN_143_1),
    ._GEN_367_0(d__GEN_367_0),
    ._GEN_247_0(d__GEN_247_0),
    ._GEN_274_0(d__GEN_274_0),
    ._GEN_460(d__GEN_460),
    ._GEN_283_0(d__GEN_283_0),
    ._GEN_388_0(d__GEN_388_0),
    ._GEN_382_0(d__GEN_382_0),
    ._GEN_268_0(d__GEN_268_0),
    ._GEN_176_1(d__GEN_176_1),
    ._GEN_346_0(d__GEN_346_0),
    ._GEN_64_1(d__GEN_64_1),
    ._GEN_340_0(d__GEN_340_0),
    ._GEN_134_1(d__GEN_134_1),
    ._GEN_149_2(d__GEN_149_2),
    ._GEN_439(d__GEN_439),
    ._GEN_262_0(d__GEN_262_0),
    ._GEN_17_1(d__GEN_17_1),
    ._GEN_361_0(d__GEN_361_0),
    ._GEN_155_1(d__GEN_155_1),
    ._GEN_170_1(d__GEN_170_1),
    ._GEN_73_1(d__GEN_73_1),
    ._GEN_128_1(d__GEN_128_1),
    ._GEN_241_0(d__GEN_241_0),
    ._GEN_445(d__GEN_445),
    ._GEN_289_0(d__GEN_289_0),
    ._GEN_131_1(d__GEN_131_1),
    ._GEN_152_2(d__GEN_152_2),
    ._GEN_421_0(d__GEN_421_0),
    ._GEN_427(d__GEN_427),
    ._GEN_454(d__GEN_454),
    ._GEN_256_0(d__GEN_256_0),
    ._GEN_110_1(d__GEN_110_1),
    ._GEN_40_1(d__GEN_40_1),
    ._GEN_5_2(d__GEN_5_2),
    ._GEN_158_1(d__GEN_158_1),
    ._GEN_271_0(d__GEN_271_0),
    ._GEN_322_0(d__GEN_322_0),
    ._GEN_334_0(d__GEN_334_0),
    ._GEN_116_1(d__GEN_116_1),
    ._GEN_235_0(d__GEN_235_0),
    ._GEN_349_0(d__GEN_349_0),
    ._GEN_147_2(d__GEN_147_2),
    ._GEN_448(d__GEN_448),
    ._GEN_442(d__GEN_442),
    ._GEN_343_0(d__GEN_343_0),
    ._GEN_355_0(d__GEN_355_0),
    ._GEN_137_1(d__GEN_137_1),
    ._GEN_370_0(d__GEN_370_0),
    ._GEN_250_0(d__GEN_250_0),
    ._GEN_463(d__GEN_463),
    ._GEN_328_0(d__GEN_328_0)
  );
  assign c_metaReset = metaReset;
  assign d_metaReset = metaReset;
  assign io_imem_req_bits_addr = d_io_imem_req_bits_addr; // @[core.scala 30:12 core.scala 31:12]
  assign io_dmem_req_valid = d_io_dmem_req_valid; // @[core.scala 34:12 core.scala 35:12]
  assign io_dmem_req_bits_addr = d_io_dmem_req_bits_addr; // @[core.scala 34:12 core.scala 35:12]
  assign io_dmem_req_bits_data = d_io_dmem_req_bits_data; // @[core.scala 34:12 core.scala 35:12]
  assign io_dmem_req_bits_fcn = d_io_dmem_req_bits_fcn; // @[core.scala 34:12 core.scala 35:12]
  assign io_dmem_req_bits_typ = d_io_dmem_req_bits_typ; // @[core.scala 34:12 core.scala 35:12]
  assign _GEN_451 = d__GEN_451;
  assign _GEN_331 = d__GEN_331;
  assign _GEN_337 = d__GEN_337;
  assign _GEN_113 = d__GEN_113_0;
  assign _GEN_111 = c__GEN_111_0;
  assign _GEN_415 = d__GEN_415;
  assign _GEN_436 = d__GEN_436;
  assign _GEN_140 = d__GEN_140_0;
  assign _GEN_71 = c__GEN_71_0;
  assign _GEN_324 = c__GEN_324_0;
  assign _GEN_219 = c__GEN_219_0;
  assign _GEN_168 = c__GEN_168_0;
  assign _GEN_98 = d__GEN_98_0;
  assign _GEN_1 = c__GEN_1_0;
  assign _GEN_352 = d__GEN_352;
  assign _GEN_423 = c__GEN_423_0;
  assign _GEN_44 = c__GEN_44_0;
  assign _GEN_125 = d__GEN_125_0;
  assign _GEN_267 = c__GEN_267_0;
  assign _GEN_126 = c__GEN_126_0;
  assign _GEN_430 = d__GEN_430;
  assign _GEN_153 = c__GEN_153_0;
  assign _GEN_225 = c__GEN_225_0;
  assign _GEN_119 = d__GEN_119_0;
  assign _GEN_88 = d__GEN_88_0;
  assign _GEN_59 = c__GEN_59_0;
  assign _GEN_252 = c__GEN_252_0;
  assign _GEN_151 = d__GEN_151_0;
  assign _GEN_147 = c__GEN_147_0;
  assign _GEN_310 = d__GEN_310;
  assign _GEN_351 = c__GEN_351_0;
  assign _GEN_210 = c__GEN_210_0;
  assign _GEN_246 = c__GEN_246_0;
  assign _GEN_104 = d__GEN_104_0;
  assign _GEN_409 = d__GEN_409;
  assign _GEN_65 = c__GEN_65_0;
  assign _GEN_253 = d__GEN_253;
  assign _GEN_132 = c__GEN_132_0;
  assign _GEN_318 = c__GEN_318_0;
  assign _GEN_316 = d__GEN_316;
  assign _GEN_92 = c__GEN_92_0;
  assign _GEN_345 = c__GEN_345_0;
  assign _GEN_231 = c__GEN_231_0;
  assign _GEN_417 = c__GEN_417_0;
  assign _GEN_244 = d__GEN_244;
  assign _GEN_50 = c__GEN_50_0;
  assign _GEN_238 = d__GEN_238;
  assign _GEN_330 = c__GEN_330_0;
  assign _GEN_86 = c__GEN_86_0;
  assign _GEN_339 = c__GEN_339_0;
  assign _GEN_101 = d__GEN_101_0;
  assign _GEN_325 = d__GEN_325;
  assign _GEN_240 = c__GEN_240_0;
  assign _GEN_234 = c__GEN_234_0;
  assign _GEN_120 = c__GEN_120_0;
  assign _GEN_169 = d__GEN_169_0;
  assign _GEN_129 = c__GEN_129_0;
  assign _GEN_433 = d__GEN_433;
  assign _GEN_333 = c__GEN_333_0;
  assign _GEN_302 = c__GEN_302_0;
  assign _GEN_313 = d__GEN_313;
  assign _GEN_228 = c__GEN_228_0;
  assign _GEN_197 = c__GEN_197_0;
  assign _GEN_91 = d__GEN_91_0;
  assign _GEN_411 = c__GEN_411_0;
  assign _GEN_11 = d__GEN_11_0;
  assign _GEN_401 = c__GEN_401_0;
  assign _GEN_47 = c__GEN_47_0;
  assign _GEN_296 = c__GEN_296_0;
  assign _GEN_304 = d__GEN_304;
  assign _GEN_294 = d__GEN_294;
  assign _GEN_74 = c__GEN_74_0;
  assign _GEN_213 = c__GEN_213_0;
  assign _GEN_303 = d__GEN_303;
  assign _GEN_107 = d__GEN_107_0;
  assign _GEN_32 = c__GEN_32_0;
  assign _GEN_0 = d__GEN_0_0;
  assign _GEN_402 = d__GEN_402;
  assign _GEN_412 = d__GEN_412;
  assign _GEN_68 = c__GEN_68_0;
  assign _GEN_135 = c__GEN_135_0;
  assign _GEN_424 = d__GEN_424;
  assign _GEN_175 = d__GEN_175_0;
  assign _GEN_319 = d__GEN_319;
  assign _GEN_288 = d__GEN_288;
  assign _GEN_56 = d__GEN_56_0;
  assign _GEN_26 = c__GEN_26_0;
  assign _GEN_418 = d__GEN_418;
  assign _GEN_122 = d__GEN_122_0;
  assign _GEN_387 = d__GEN_387;
  assign _GEN_53 = c__GEN_53_0;
  assign _GEN_141 = c__GEN_141_0;
  assign _GEN_327 = c__GEN_327_0;
  assign _GEN_72 = d__GEN_72_0;
  assign _GEN_395 = c__GEN_395_0;
  assign _GEN_249 = c__GEN_249_0;
  assign _GEN_114 = c__GEN_114_0;
  assign _GEN_312 = c__GEN_312_0;
  assign _GEN_203 = c__GEN_203_0;
  assign _GEN_75 = d__GEN_75_0;
  assign _GEN_85 = d__GEN_85_0;
  assign _GEN_20 = c__GEN_20_0;
  assign _GEN_178 = d__GEN_178_0;
  assign _GEN_15 = c__GEN_15_0;
  assign _GEN_157 = d__GEN_157_0;
  assign _GEN_462 = d__GEN_462;
  assign _GEN_69 = d__GEN_69_0;
  assign _GEN_216 = c__GEN_216_0;
  assign _GEN_206 = c__GEN_206_0;
  assign _GEN_375 = d__GEN_375;
  assign _GEN_151_0 = d__GEN_151_1;
  assign _GEN_420 = c__GEN_420_0;
  assign _GEN_123 = c__GEN_123_0;
  assign _GEN_315 = c__GEN_315_0;
  assign _GEN_284 = c__GEN_284_0;
  assign _GEN_179 = c__GEN_179_0;
  assign _GEN_33 = d__GEN_33_0;
  assign _GEN_222 = c__GEN_222_0;
  assign _GEN_377 = c__GEN_377_0;
  assign _GEN_191 = c__GEN_191_0;
  assign _GEN_290 = c__GEN_290_0;
  assign _GEN_404 = c__GEN_404_0;
  assign _GEN_390 = d__GEN_390;
  assign _GEN_56_0 = c__GEN_56_1;
  assign _GEN_305 = c__GEN_305_0;
  assign _GEN_299 = c__GEN_299_0;
  assign _GEN_185 = c__GEN_185_0;
  assign _GEN_307 = d__GEN_307;
  assign _GEN_297 = d__GEN_297;
  assign _GEN_398 = c__GEN_398_0;
  assign _GEN_406 = d__GEN_406;
  assign _GEN_41 = c__GEN_41_0;
  assign _GEN_321 = c__GEN_321_0;
  assign _GEN_270 = d__GEN_270;
  assign _GEN_95 = d__GEN_95_0;
  assign _GEN_45 = d__GEN_45_0;
  assign _GEN_414 = c__GEN_414_0;
  assign _GEN_383 = c__GEN_383_0;
  assign _GEN_369 = d__GEN_369;
  assign _GEN_35 = c__GEN_35_0;
  assign _GEN_29 = c__GEN_29_0;
  assign _GEN_278 = c__GEN_278_0;
  assign _GEN_117 = c__GEN_117_0;
  assign _GEN_396 = d__GEN_396;
  assign _GEN_172 = d__GEN_172_0;
  assign _GEN_276 = d__GEN_276;
  assign _GEN_291 = d__GEN_291;
  assign _GEN_365 = c__GEN_365_0;
  assign _GEN_359 = c__GEN_359_0;
  assign _GEN_258 = d__GEN_258;
  assign _GEN_372 = d__GEN_372;
  assign _GEN_38 = c__GEN_38_0;
  assign _GEN_252_0 = d__GEN_252_0;
  assign _GEN_167 = c__GEN_167_0;
  assign _GEN_166 = d__GEN_166_0;
  assign _GEN_285 = d__GEN_285;
  assign _GEN_42 = d__GEN_42_0;
  assign _GEN_350 = c__GEN_350_0;
  assign _GEN_106 = c__GEN_106_0;
  assign _GEN_384 = d__GEN_384;
  assign _GEN_18 = c__GEN_18_0;
  assign _GEN_378 = d__GEN_378;
  assign _GEN_393 = d__GEN_393;
  assign _GEN_273 = d__GEN_273;
  assign _GEN_293 = c__GEN_293_0;
  assign _GEN_456 = d__GEN_456;
  assign _GEN_371 = c__GEN_371_0;
  assign _GEN_80 = d__GEN_80_0;
  assign _GEN_351_0 = d__GEN_351_0;
  assign _GEN_251 = c__GEN_251_0;
  assign _GEN_209 = c__GEN_209_0;
  assign _GEN_139 = d__GEN_139_0;
  assign _GEN_145 = d__GEN_145_0;
  assign _GEN_450 = d__GEN_450;
  assign _GEN_308 = c__GEN_308_0;
  assign _GEN_173 = c__GEN_173_0;
  assign _GEN_53_0 = d__GEN_53_1;
  assign _GEN_357 = d__GEN_357;
  assign _GEN_200 = c__GEN_200_0;
  assign _GEN_386 = c__GEN_386_0;
  assign _GEN_272 = c__GEN_272_0;
  assign _GEN_160 = d__GEN_160_0;
  assign _GEN_91_0 = c__GEN_91_1;
  assign _GEN_279 = d__GEN_279;
  assign _GEN_194 = c__GEN_194_0;
  assign _GEN_188 = c__GEN_188_0;
  assign _GEN_133 = d__GEN_133_0;
  assign _GEN_392 = c__GEN_392_0;
  assign _GEN_23 = c__GEN_23_0;
  assign _GEN_407 = c__GEN_407_0;
  assign _GEN_287 = c__GEN_287_0;
  assign _GEN_266 = c__GEN_266_0;
  assign _GEN_399 = d__GEN_399;
  assign _GEN_264 = d__GEN_264;
  assign _GEN_300 = d__GEN_300;
  assign _GEN_374 = c__GEN_374_0;
  assign _GEN_233 = c__GEN_233_0;
  assign _GEN_127 = d__GEN_127_0;
  assign _GEN_269 = c__GEN_269_0;
  assign _GEN_432 = d__GEN_432;
  assign _GEN_381 = d__GEN_381;
  assign _GEN_260 = c__GEN_260_0;
  assign _GEN_161 = c__GEN_161_0;
  assign _GEN_155 = c__GEN_155_0;
  assign _GEN_339_0 = d__GEN_339_0;
  assign _GEN_368 = c__GEN_368_0;
  assign _GEN_254 = c__GEN_254_0;
  assign _GEN_281 = c__GEN_281_0;
  assign _GEN_73 = c__GEN_73_0;
  assign _GEN_261 = d__GEN_261;
  assign _GEN_353 = c__GEN_353_0;
  assign _GEN_332 = c__GEN_332_0;
  assign _GEN_88_0 = c__GEN_88_1;
  assign _GEN_176 = c__GEN_176_0;
  assign _GEN_16 = d__GEN_16_0;
  assign _GEN_380 = c__GEN_380_0;
  assign _GEN_360 = d__GEN_360;
  assign _GEN_389 = c__GEN_389_0;
  assign _GEN_163 = d__GEN_163_0;
  assign _GEN_246_0 = d__GEN_246_0;
  assign _GEN_438 = d__GEN_438;
  assign _GEN_94 = c__GEN_94_0;
  assign _GEN_282 = d__GEN_282;
  assign _GEN_347 = c__GEN_347_0;
  assign _GEN_109 = c__GEN_109_0;
  assign _GEN_182 = c__GEN_182_0;
  assign _GEN_345_0 = d__GEN_345_0;
  assign _GEN_121 = d__GEN_121_0;
  assign _GEN_240_0 = d__GEN_240_0;
  assign _GEN_9 = c__GEN_9_0;
  assign _GEN_148 = d__GEN_148_0;
  assign _GEN_154 = d__GEN_154_0;
  assign _GEN_444 = d__GEN_444;
  assign _GEN_149 = c__GEN_149_0;
  assign _GEN_267_0 = d__GEN_267_0;
  assign _GEN_459 = d__GEN_459;
  assign _GEN_453 = d__GEN_453;
  assign _GEN_248 = c__GEN_248_0;
  assign _GEN_366 = d__GEN_366;
  assign _GEN_7 = d__GEN_7_0;
  assign _GEN_142 = d__GEN_142_0;
  assign _GEN_275 = c__GEN_275_0;
  assign _GEN_140_0 = c__GEN_140_1;
  assign _GEN_324_0 = d__GEN_324_0;
  assign _GEN_100 = c__GEN_100_0;
  assign _GEN_333_0 = d__GEN_333_0;
  assign _GEN_362 = c__GEN_362_0;
  assign _GEN_413 = c__GEN_413_0;
  assign _GEN_342 = d__GEN_342;
  assign _GEN_405 = d__GEN_405;
  assign _GEN_420_0 = d__GEN_420_0;
  assign _GEN_306 = d__GEN_306;
  assign _GEN_76 = c__GEN_76_0;
  assign _GEN_164 = c__GEN_164_0;
  assign _GEN_109_0 = d__GEN_109_1;
  assign _GEN_103 = d__GEN_103_0;
  assign _GEN_3 = d__GEN_3_0;
  assign _GEN_242 = c__GEN_242_0;
  assign _GEN_136 = d__GEN_136_0;
  assign _GEN_426 = d__GEN_426;
  assign _GEN_137 = c__GEN_137_0;
  assign _GEN_441 = d__GEN_441;
  assign _GEN_341 = c__GEN_341_0;
  assign _GEN_94_0 = d__GEN_94_1;
  assign _GEN_348 = d__GEN_348;
  assign _GEN_263 = c__GEN_263_0;
  assign _GEN_257 = c__GEN_257_0;
  assign _GEN_122_0 = c__GEN_122_1;
  assign _GEN_143 = c__GEN_143_0;
  assign _GEN_255 = d__GEN_255;
  assign _GEN_82 = c__GEN_82_0;
  assign _GEN_170 = c__GEN_170_0;
  assign _GEN_356 = c__GEN_356_0;
  assign _GEN_221 = c__GEN_221_0;
  assign _GEN_215 = c__GEN_215_0;
  assign _GEN_115 = d__GEN_115_0;
  assign _GEN_146 = d__GEN_146_0;
  assign _GEN_363 = d__GEN_363;
  assign _GEN_320 = c__GEN_320_0;
  assign _GEN_314 = c__GEN_314_0;
  assign _GEN_329 = c__GEN_329_0;
  assign _GEN_321_0 = d__GEN_321_0;
  assign _GEN_327_0 = d__GEN_327_0;
  assign _GEN_103_0 = c__GEN_103_1;
  assign _GEN_97 = c__GEN_97_0;
  assign _GEN_236 = c__GEN_236_0;
  assign _GEN_354 = d__GEN_354;
  assign _GEN_234_0 = d__GEN_234_0;
  assign _GEN_130 = d__GEN_130_0;
  assign _GEN_61 = c__GEN_61_0;
  assign _GEN_55 = c__GEN_55_0;
  assign _GEN_249_0 = d__GEN_249_0;
  assign _GEN_335 = c__GEN_335_0;
  assign _GEN_243 = d__GEN_243;
  assign _GEN_447 = d__GEN_447;
  assign _GEN_158 = c__GEN_158_0;
  assign _GEN_330_0 = d__GEN_330_0;
  assign _GEN_422 = c__GEN_422_0;
  assign _GEN_245 = c__GEN_245_0;
  assign _GEN_37 = c__GEN_37_0;
  assign _GEN_125_0 = c__GEN_125_1;
  assign _GEN_429 = d__GEN_429;
  assign _GEN_70 = c__GEN_70_0;
  assign _GEN_64 = c__GEN_64_0;
  assign _GEN_344 = c__GEN_344_0;
  assign _GEN_338 = c__GEN_338_0;
  assign _GEN_293_0 = d__GEN_293_0;
  assign _GEN_87 = d__GEN_87_0;
  assign _GEN_416 = c__GEN_416_0;
  assign _GEN_406_0 = c__GEN_406_1;
  assign _GEN_58 = c__GEN_58_0;
  assign _GEN_414_0 = d__GEN_414_0;
  assign _GEN_309 = d__GEN_309;
  assign _GEN_85_0 = c__GEN_85_1;
  assign _GEN_299_0 = d__GEN_299_0;
  assign _GEN_336 = d__GEN_336;
  assign _GEN_408 = d__GEN_408;
  assign _GEN_112 = d__GEN_112_0;
  assign _GEN_43 = c__GEN_43_0;
  assign _GEN_150 = d__GEN_150_0;
  assign _GEN_131 = c__GEN_131_0;
  assign _GEN_435 = d__GEN_435;
  assign _GEN_230 = c__GEN_230_0;
  assign _GEN_97_0 = d__GEN_97_1;
  assign _GEN_124 = d__GEN_124_0;
  assign _GEN_239 = c__GEN_239_0;
  assign _GEN_118 = d__GEN_118_0;
  assign _GEN_392_0 = d__GEN_392_0;
  assign _GEN_398_0 = d__GEN_398_0;
  assign _GEN_423_0 = d__GEN_423_0;
  assign _GEN_237 = d__GEN_237;
  assign _GEN_152 = c__GEN_152_0;
  assign _GEN_307_0 = c__GEN_307_1;
  assign _GEN_146_0 = c__GEN_146_1;
  assign _GEN_315_0 = d__GEN_315_0;
  assign _GEN_79 = d__GEN_79_0;
  assign _GEN_224 = c__GEN_224_0;
  assign _GEN_110 = c__GEN_110_0;
  assign _GEN_119_0 = c__GEN_119_1;
  assign _GEN_323 = c__GEN_323_0;
  assign _GEN_317 = c__GEN_317_0;
  assign _GEN_79_0 = c__GEN_79_1;
  assign _GEN_218 = c__GEN_218_0;
  assign _GEN_208 = c__GEN_208_0;
  assign _GEN_1_1 = d__GEN_1_2;
  assign _GEN_196 = c__GEN_196_0;
  assign _GEN_90 = d__GEN_90_0;
  assign _GEN_31 = c__GEN_31_0;
  assign _GEN_400 = c__GEN_400_0;
  assign _GEN_113_0 = c__GEN_113_1;
  assign _GEN_162 = d__GEN_162_0;
  assign _GEN_212 = c__GEN_212_0;
  assign _GEN_302_0 = d__GEN_302_0;
  assign _GEN_181 = c__GEN_181_0;
  assign _GEN_106_0 = d__GEN_106_1;
  assign _GEN_227 = c__GEN_227_0;
  assign _GEN_71_0 = d__GEN_71_1;
  assign _GEN_380_0 = d__GEN_380_0;
  assign _GEN_425 = c__GEN_425_0;
  assign _GEN_280 = c__GEN_280_0;
  assign _GEN_46 = c__GEN_46_0;
  assign _GEN_174 = d__GEN_174_0;
  assign _GEN_134 = c__GEN_134_0;
  assign _GEN_289 = c__GEN_289_0;
  assign _GEN_318_0 = d__GEN_318_0;
  assign _GEN_287_0 = d__GEN_287_0;
  assign _GEN_202 = c__GEN_202_0;
  assign _GEN_419 = c__GEN_419_0;
  assign _GEN_388 = c__GEN_388_0;
  assign _GEN_410 = c__GEN_410_0;
  assign _GEN_386_0 = d__GEN_386_0;
  assign _GEN_52 = c__GEN_52_0;
  assign _GEN_311 = c__GEN_311_0;
  assign _GEN_301 = c__GEN_301_0;
  assign _GEN_295 = c__GEN_295_0;
  assign _GEN_67 = c__GEN_67_0;
  assign _GEN_281_0 = d__GEN_281_0;
  assign _GEN_312_0 = d__GEN_312_0;
  assign _GEN_25 = c__GEN_25_0;
  assign _GEN_409_0 = c__GEN_409_1;
  assign _GEN_417_0 = d__GEN_417_0;
  assign _GEN_411_0 = d__GEN_411_0;
  assign _GEN_326 = c__GEN_326_0;
  assign _GEN_55_0 = d__GEN_55_1;
  assign _GEN_100_0 = d__GEN_100_1;
  assign _GEN_394 = c__GEN_394_0;
  assign _GEN_168_0 = d__GEN_168_1;
  assign _GEN_128 = c__GEN_128_0;
  assign _GEN_401_0 = d__GEN_401_0;
  assign _GEN_44_0 = d__GEN_44_1;
  assign _GEN_376 = c__GEN_376_0;
  assign _GEN_74_0 = d__GEN_74_1;
  assign _GEN_374_0 = d__GEN_374_0;
  assign _GEN_40 = c__GEN_40_0;
  assign _GEN_368_0 = d__GEN_368_0;
  assign _GEN_34 = c__GEN_34_0;
  assign _GEN_383_0 = d__GEN_383_0;
  assign _GEN_49 = c__GEN_49_0;
  assign _GEN_263_0 = d__GEN_263_0;
  assign _GEN_177 = d__GEN_177_0;
  assign _GEN_171 = d__GEN_171_0;
  assign _GEN_446 = d__GEN_446;
  assign _GEN_102 = c__GEN_102_0;
  assign _GEN_290_0 = d__GEN_290_0;
  assign _GEN_190 = c__GEN_190_0;
  assign _GEN_83 = d__GEN_83_0;
  assign _GEN_205 = c__GEN_205_0;
  assign _GEN_135_0 = d__GEN_135_1;
  assign _GEN_389_0 = d__GEN_389_0;
  assign _GEN_93 = d__GEN_93_0;
  assign _GEN_254_0 = d__GEN_254_0;
  assign _GEN_298 = c__GEN_298_0;
  assign _GEN_163_0 = c__GEN_163_1;
  assign _GEN_21 = d__GEN_21_0;
  assign _GEN_461 = d__GEN_461;
  assign _GEN_362_0 = d__GEN_362_0;
  assign _GEN_14 = c__GEN_14_0;
  assign _GEN_116 = c__GEN_116_0;
  assign _GEN_156 = d__GEN_156_0;
  assign _GEN_150_0 = d__GEN_150_1;
  assign _GEN_283 = c__GEN_283_0;
  assign _GEN_184 = c__GEN_184_0;
  assign _GEN_178_0 = c__GEN_178_1;
  assign _GEN_68_0 = d__GEN_68_1;
  assign _GEN_296_0 = d__GEN_296_0;
  assign _GEN_382 = c__GEN_382_0;
  assign _GEN_397 = c__GEN_397_0;
  assign _GEN_277 = c__GEN_277_0;
  assign _GEN_395_0 = d__GEN_395_0;
  assign _GEN_304_0 = c__GEN_304_1;
  assign _GEN_199 = c__GEN_199_0;
  assign _GEN_403 = c__GEN_403_0;
  assign _GEN_262 = c__GEN_262_0;
  assign _GEN_28 = c__GEN_28_0;
  assign _GEN_275_0 = d__GEN_275_0;
  assign _GEN_269_0 = d__GEN_269_0;
  assign _GEN_361 = c__GEN_361_0;
  assign _GEN_96 = c__GEN_96_0;
  assign _GEN_278_0 = d__GEN_278_0;
  assign _GEN_193 = c__GEN_193_0;
  assign _GEN_379 = c__GEN_379_0;
  assign _GEN_244_0 = c__GEN_244_1;
  assign _GEN_138 = d__GEN_138_0;
  assign _GEN_271 = c__GEN_271_0;
  assign _GEN_251_0 = d__GEN_251_0;
  assign _GEN_151_1 = c__GEN_151_2;
  assign _GEN_166_0 = c__GEN_166_1;
  assign _GEN_455 = d__GEN_455;
  assign _GEN_370 = c__GEN_370_0;
  assign _GEN_364 = c__GEN_364_0;
  assign _GEN_259 = c__GEN_259_0;
  assign _GEN_377_0 = d__GEN_377_0;
  assign _GEN_153_0 = d__GEN_153_1;
  assign _GEN_292 = c__GEN_292_0;
  assign _GEN_84 = c__GEN_84_0;
  assign _GEN_78 = c__GEN_78_0;
  assign _GEN_272_0 = d__GEN_272_0;
  assign _GEN_47_0 = d__GEN_47_1;
  assign _GEN_335_0 = d__GEN_335_0;
  assign _GEN_41_0 = d__GEN_41_1;
  assign _GEN_385 = c__GEN_385_0;
  assign _GEN_250 = c__GEN_250_0;
  assign _GEN_434 = d__GEN_434;
  assign _GEN_257_0 = d__GEN_257_0;
  assign _GEN_343 = c__GEN_343_0;
  assign _GEN_443 = d__GEN_443;
  assign _GEN_105 = c__GEN_105_0;
  assign _GEN_99 = c__GEN_99_0;
  assign _GEN_358 = c__GEN_358_0;
  assign _GEN_356_0 = d__GEN_356_0;
  assign _GEN_350_0 = d__GEN_350_0;
  assign _GEN_132_0 = d__GEN_132_1;
  assign _GEN_22 = c__GEN_22_0;
  assign _GEN_144 = d__GEN_144_0;
  assign _GEN_265 = c__GEN_265_0;
  assign _GEN_17 = c__GEN_17_0;
  assign _GEN_159 = d__GEN_159_0;
  assign _GEN_428 = d__GEN_428;
  assign _GEN_449 = d__GEN_449;
  assign _GEN_90_0 = c__GEN_90_1;
  assign _GEN_172_0 = c__GEN_172_1;
  assign _GEN_187 = c__GEN_187_0;
  assign _GEN_117_0 = d__GEN_117_1;
  assign _GEN_236_0 = d__GEN_236_0;
  assign _GEN_371_0 = d__GEN_371_0;
  assign _GEN_391 = c__GEN_391_0;
  assign _GEN_165 = d__GEN_165_0;
  assign _GEN_286 = c__GEN_286_0;
  assign _GEN_145_0 = c__GEN_145_1;
  assign _GEN_284_0 = d__GEN_284_0;
  assign _GEN_232 = c__GEN_232_0;
  assign _GEN_147_0 = d__GEN_147_1;
  assign _GEN_416_0 = d__GEN_416_0;
  assign _GEN_274 = c__GEN_274_0;
  assign _GEN_260_0 = d__GEN_260_0;
  assign _GEN_175_0 = c__GEN_175_1;
  assign _GEN_105_0 = d__GEN_105_1;
  assign _GEN_169_0 = c__GEN_169_1;
  assign _GEN_338_0 = d__GEN_338_0;
  assign _GEN_247 = c__GEN_247_0;
  assign _GEN_133_0 = c__GEN_133_1;
  assign _GEN_141_0 = d__GEN_141_1;
  assign _GEN_160_0 = c__GEN_160_1;
  assign _GEN_346 = c__GEN_346_0;
  assign _GEN_99_0 = d__GEN_99_1;
  assign _GEN_344_0 = d__GEN_344_0;
  assign _GEN_373 = c__GEN_373_0;
  assign _GEN_424_0 = c__GEN_424_1;
  assign _GEN_239_0 = d__GEN_239_0;
  assign _GEN_353_0 = d__GEN_353_0;
  assign _GEN_268 = c__GEN_268_0;
  assign _GEN_127_0 = c__GEN_127_1;
  assign _GEN_8 = c__GEN_8_0;
  assign _GEN_266_0 = d__GEN_266_0;
  assign _GEN_331_0 = c__GEN_331_1;
  assign _GEN_452 = d__GEN_452;
  assign _GEN_93_0 = c__GEN_93_1;
  assign _GEN_87_0 = c__GEN_87_1;
  assign _GEN_367 = c__GEN_367_0;
  assign _GEN_226 = c__GEN_226_0;
  assign _GEN_120_0 = d__GEN_120_1;
  assign _GEN_365_0 = d__GEN_365_0;
  assign _GEN_6 = d__GEN_6_0;
  assign _GEN_410_0 = d__GEN_410_0;
  assign _GEN_253_0 = c__GEN_253_1;
  assign _GEN_152_0 = d__GEN_152_1;
  assign _GEN_325_0 = c__GEN_325_1;
  assign _GEN_148_0 = c__GEN_148_1;
  assign _GEN_437 = d__GEN_437;
  assign _GEN_352_0 = c__GEN_352_1;
  assign _GEN_332_0 = d__GEN_332_0;
  assign _GEN_108 = c__GEN_108_0;
  assign _GEN_126_0 = d__GEN_126_1;
  assign _GEN_245_0 = d__GEN_245_0;
  assign _GEN_359_0 = d__GEN_359_0;
  assign _GEN_431 = d__GEN_431;
  assign _GEN_72_0 = c__GEN_72_1;
  assign _GEN_66 = c__GEN_66_0;
  assign _GEN_154_0 = c__GEN_154_1;
  assign _GEN_458 = d__GEN_458;
  assign _GEN_317_0 = d__GEN_317_0;
  assign _GEN_326_0 = d__GEN_326_0;
  assign _GEN_241 = c__GEN_241_0;
  assign _GEN_341_0 = d__GEN_341_0;
  assign _GEN_402_0 = c__GEN_402_1;
  assign _GEN_1_2 = d__GEN_1_3;
  assign _GEN_48 = c__GEN_48_0;
  assign _GEN_394_0 = d__GEN_394_0;
  assign _GEN_60 = c__GEN_60_0;
  assign _GEN_248_0 = d__GEN_248_0;
  assign _GEN_75_0 = c__GEN_75_1;
  assign _GEN_349 = c__GEN_349_0;
  assign _GEN_214 = c__GEN_214_0;
  assign _GEN_347_0 = d__GEN_347_0;
  assign _GEN_412_0 = c__GEN_412_1;
  assign _GEN_92_0 = d__GEN_92_1;
  assign _GEN_102_0 = d__GEN_102_1;
  assign _GEN_256 = c__GEN_256_0;
  assign _GEN_121_0 = c__GEN_121_1;
  assign _GEN_425_0 = d__GEN_425_0;
  assign _GEN_305_0 = d__GEN_305_0;
  assign _GEN_419_0 = d__GEN_419_0;
  assign _GEN_81 = c__GEN_81_0;
  assign _GEN_320_0 = d__GEN_320_0;
  assign _GEN_108_0 = d__GEN_108_1;
  assign _GEN_114_0 = d__GEN_114_1;
  assign _GEN_123_0 = d__GEN_123_1;
  assign _GEN_413_0 = d__GEN_413_0;
  assign _GEN_54 = c__GEN_54_0;
  assign _GEN_136_0 = c__GEN_136_1;
  assign _GEN_142_0 = c__GEN_142_1;
  assign _GEN_440 = d__GEN_440;
  assign _GEN_295_0 = d__GEN_295_0;
  assign _GEN_340 = c__GEN_340_0;
  assign _GEN_355 = c__GEN_355_0;
  assign _GEN_235 = c__GEN_235_0;
  assign _GEN_129_0 = d__GEN_129_1;
  assign _GEN_404_0 = d__GEN_404_0;
  assign _GEN_403_0 = d__GEN_403_0;
  assign _GEN_313_0 = c__GEN_313_1;
  assign _GEN_242_0 = d__GEN_242_0;
  assign _GEN_69_0 = c__GEN_69_1;
  assign _GEN_157_0 = c__GEN_157_1;
  assign _GEN_220 = c__GEN_220_0;
  assign _GEN_229 = c__GEN_229_0;
  assign _GEN_115_0 = c__GEN_115_1;
  assign _GEN_15_0 = d__GEN_15_1;
  assign _GEN_334 = c__GEN_334_0;
  assign _GEN_328 = c__GEN_328_0;
  assign _GEN_96_0 = d__GEN_96_1;
  assign _GEN_86_0 = d__GEN_86_1;
  assign _GEN_36 = c__GEN_36_0;
  assign _GEN_405_0 = c__GEN_405_1;
  assign _GEN_415_0 = c__GEN_415_1;
  assign _GEN_164_0 = d__GEN_164_1;
  assign _GEN_124_0 = c__GEN_124_1;
  assign _GEN_322 = c__GEN_322_0;
  assign _GEN_308_0 = d__GEN_308_0;
  assign _GEN_337_0 = c__GEN_337_1;
  assign _GEN_223 = c__GEN_223_0;
  assign _GEN_217 = c__GEN_217_0;
  assign _GEN_192 = c__GEN_192_0;
  assign _GEN_390_0 = c__GEN_390_1;
  assign _GEN_42_0 = c__GEN_42_1;
  assign _GEN_149_0 = d__GEN_149_1;
  assign _GEN_291_0 = c__GEN_291_1;
  assign _GEN_139_0 = c__GEN_139_1;
  assign _GEN_329_0 = d__GEN_329_0;
  assign _GEN_292_0 = d__GEN_292_0;
  assign _GEN_298_0 = d__GEN_298_0;
  assign _GEN_207 = c__GEN_207_0;
  assign _GEN_399_0 = c__GEN_399_1;
  assign _GEN_421 = c__GEN_421_0;
  assign _GEN_63 = c__GEN_63_0;
  assign _GEN_391_0 = d__GEN_391_0;
  assign _GEN_316_0 = c__GEN_316_1;
  assign _GEN_306_0 = c__GEN_306_1;
  assign _GEN_314_0 = d__GEN_314_0;
  assign _GEN_21_0 = c__GEN_21_1;
  assign _GEN_323_0 = d__GEN_323_0;
  assign _GEN_384_0 = c__GEN_384_1;
  assign _GEN_118_0 = c__GEN_118_1;
  assign _GEN_376_0 = d__GEN_376_0;
  assign _GEN_422_0 = d__GEN_422_0;
  assign _GEN_277_0 = d__GEN_277_0;
  assign _GEN_57 = c__GEN_57_0;
  assign _GEN_130_0 = c__GEN_130_1;
  assign _GEN_46_0 = d__GEN_46_1;
  assign _GEN_111_0 = d__GEN_111_1;
  assign _GEN_78_0 = d__GEN_78_1;
  assign _GEN_238_0 = c__GEN_238_1;
  assign _GEN_407_0 = d__GEN_407_0;
  assign _GEN_179_0 = d__GEN_179_1;
  assign _GEN_397_0 = d__GEN_397_0;
  assign _GEN_173_0 = d__GEN_173_1;
  assign _GEN_70_0 = d__GEN_70_1;
  assign _GEN_379_0 = d__GEN_379_0;
  assign _GEN_82_0 = d__GEN_82_1;
  assign _GEN_373_0 = d__GEN_373_0;
  assign _GEN_45_0 = c__GEN_45_1;
  assign _GEN_54_0 = d__GEN_54_1;
  assign _GEN_201 = c__GEN_201_0;
  assign _GEN_195 = c__GEN_195_0;
  assign _GEN_364_0 = d__GEN_364_0;
  assign _GEN_259_0 = d__GEN_259_0;
  assign _GEN_167_0 = d__GEN_167_1;
  assign _GEN_309_0 = c__GEN_309_1;
  assign _GEN_43_0 = d__GEN_43_1;
  assign _GEN_372_0 = c__GEN_372_1;
  assign _GEN_19 = c__GEN_19_0;
  assign _GEN_161_0 = d__GEN_161_1;
  assign _GEN_51 = c__GEN_51_0;
  assign _GEN_265_0 = d__GEN_265_0;
  assign _GEN_294_0 = c__GEN_294_1;
  assign _GEN_180 = c__GEN_180_0;
  assign _GEN_189 = c__GEN_189_0;
  assign _GEN_211 = c__GEN_211_0;
  assign _GEN_301_0 = d__GEN_301_0;
  assign _GEN_393_0 = c__GEN_393_1;
  assign _GEN_387_0 = c__GEN_387_1;
  assign _GEN_39 = c__GEN_39_0;
  assign _GEN_146_1 = d__GEN_146_2;
  assign _GEN_288_0 = c__GEN_288_1;
  assign _GEN_310_0 = c__GEN_310_1;
  assign _GEN_300_0 = c__GEN_300_1;
  assign _GEN_286_0 = d__GEN_286_0;
  assign _GEN_400_0 = d__GEN_400_0;
  assign _GEN_319_0 = c__GEN_319_1;
  assign _GEN_107_0 = c__GEN_107_1;
  assign _GEN_174_0 = c__GEN_174_1;
  assign _GEN_89 = d__GEN_89_0;
  assign _GEN_358_0 = d__GEN_358_0;
  assign _GEN_30 = c__GEN_30_0;
  assign _GEN_24 = c__GEN_24_0;
  assign _GEN_408_0 = c__GEN_408_1;
  assign _GEN_418_0 = c__GEN_418_1;
  assign _GEN_273_0 = c__GEN_273_1;
  assign _GEN_5_0 = c__GEN_5_1;
  assign _GEN_112_0 = c__GEN_112_1;
  assign _GEN_385_0 = d__GEN_385_0;
  assign _GEN_457 = d__GEN_457;
  assign _GEN_311_0 = d__GEN_311_0;
  assign _GEN_280_0 = d__GEN_280_0;
  assign _GEN_366_0 = c__GEN_366_1;
  assign _GEN_360_0 = c__GEN_360_1;
  assign _GEN_354_0 = c__GEN_354_1;
  assign _GEN_143_0 = d__GEN_143_1;
  assign _GEN_367_0 = d__GEN_367_0;
  assign _GEN_33_0 = c__GEN_33_1;
  assign _GEN_247_0 = d__GEN_247_0;
  assign _GEN_276_0 = c__GEN_276_1;
  assign _GEN_348_0 = c__GEN_348_1;
  assign _GEN_274_0 = d__GEN_274_0;
  assign _GEN_460 = d__GEN_460;
  assign _GEN_101_0 = c__GEN_101_1;
  assign _GEN_375_0 = c__GEN_375_1;
  assign _GEN_283_0 = d__GEN_283_0;
  assign _GEN_27 = c__GEN_27_0;
  assign _GEN_13 = c__GEN_13_0;
  assign _GEN_388_0 = d__GEN_388_0;
  assign _GEN_382_0 = d__GEN_382_0;
  assign _GEN_268_0 = d__GEN_268_0;
  assign _GEN_297_0 = c__GEN_297_1;
  assign _GEN_89_0 = c__GEN_89_1;
  assign _GEN_176_0 = d__GEN_176_1;
  assign _GEN_177_0 = c__GEN_177_1;
  assign _GEN_346_0 = d__GEN_346_0;
  assign _GEN_64_0 = d__GEN_64_1;
  assign _GEN_340_0 = d__GEN_340_0;
  assign _GEN_255_0 = c__GEN_255_1;
  assign _GEN_204 = c__GEN_204_0;
  assign _GEN_134_0 = d__GEN_134_1;
  assign _GEN_149_1 = d__GEN_149_2;
  assign _GEN_439 = d__GEN_439;
  assign _GEN_80_0 = c__GEN_80_1;
  assign _GEN_262_0 = d__GEN_262_0;
  assign _GEN_303_0 = c__GEN_303_1;
  assign _GEN_162_0 = c__GEN_162_1;
  assign _GEN_17_0 = d__GEN_17_1;
  assign _GEN_198 = c__GEN_198_0;
  assign _GEN_361_0 = d__GEN_361_0;
  assign _GEN_381_0 = c__GEN_381_1;
  assign _GEN_261_0 = c__GEN_261_1;
  assign _GEN_155_0 = d__GEN_155_1;
  assign _GEN_156_0 = c__GEN_156_1;
  assign _GEN_170_0 = d__GEN_170_1;
  assign _GEN_95_0 = c__GEN_95_1;
  assign _GEN_183 = c__GEN_183_0;
  assign _GEN_369_0 = c__GEN_369_1;
  assign _GEN_73_0 = d__GEN_73_1;
  assign _GEN_128_0 = d__GEN_128_1;
  assign _GEN_241_0 = d__GEN_241_0;
  assign _GEN_282_0 = c__GEN_282_1;
  assign _GEN_396_0 = c__GEN_396_1;
  assign _GEN_445 = d__GEN_445;
  assign _GEN_289_0 = d__GEN_289_0;
  assign _GEN_378_0 = c__GEN_378_1;
  assign _GEN_186 = c__GEN_186_0;
  assign _GEN_131_0 = d__GEN_131_1;
  assign _GEN_152_1 = d__GEN_152_2;
  assign _GEN_421_0 = d__GEN_421_0;
  assign _GEN_427 = d__GEN_427;
  assign _GEN_62 = c__GEN_62_0;
  assign _GEN_285_0 = c__GEN_285_1;
  assign _GEN_336_0 = c__GEN_336_1;
  assign _GEN_144_0 = c__GEN_144_1;
  assign _GEN_150_1 = c__GEN_150_2;
  assign _GEN_454 = d__GEN_454;
  assign _GEN_363_0 = c__GEN_363_1;
  assign _GEN_243_0 = c__GEN_243_1;
  assign _GEN_258_0 = c__GEN_258_1;
  assign _GEN_138_0 = c__GEN_138_1;
  assign _GEN_256_0 = d__GEN_256_0;
  assign _GEN_171_0 = c__GEN_171_1;
  assign _GEN_357_0 = c__GEN_357_1;
  assign _GEN_165_0 = c__GEN_165_1;
  assign _GEN_110_0 = d__GEN_110_1;
  assign _GEN_40_0 = d__GEN_40_1;
  assign _GEN_264_0 = c__GEN_264_1;
  assign _GEN_5_1 = d__GEN_5_2;
  assign _GEN_158_0 = d__GEN_158_1;
  assign _GEN_16_0 = c__GEN_16_1;
  assign _GEN_271_0 = d__GEN_271_0;
  assign _GEN_342_0 = c__GEN_342_1;
  assign _GEN_322_0 = d__GEN_322_0;
  assign _GEN_98_0 = c__GEN_98_1;
  assign _GEN_237_0 = c__GEN_237_1;
  assign _GEN_334_0 = d__GEN_334_0;
  assign _GEN_116_0 = d__GEN_116_1;
  assign _GEN_235_0 = d__GEN_235_0;
  assign _GEN_349_0 = d__GEN_349_0;
  assign _GEN_147_1 = d__GEN_147_2;
  assign _GEN_448 = d__GEN_448;
  assign _GEN_442 = d__GEN_442;
  assign _GEN_83_0 = c__GEN_83_1;
  assign _GEN_343_0 = d__GEN_343_0;
  assign _GEN_355_0 = d__GEN_355_0;
  assign _GEN_137_0 = d__GEN_137_1;
  assign _GEN_370_0 = d__GEN_370_0;
  assign _GEN_250_0 = d__GEN_250_0;
  assign _GEN_77 = c__GEN_77_0;
  assign _GEN_270_0 = c__GEN_270_1;
  assign _GEN_279_0 = c__GEN_279_1;
  assign _GEN_159_0 = c__GEN_159_1;
  assign _GEN_463 = d__GEN_463;
  assign _GEN_328_0 = d__GEN_328_0;
  assign _GEN_104_0 = c__GEN_104_1;
  assign c_clock = clock;
  assign c_reset = reset;
  assign c_io_imem_resp_valid = io_imem_resp_valid; // @[core.scala 30:12]
  assign c_io_dmem_resp_valid = io_dmem_resp_valid; // @[core.scala 34:12]
  assign c_io_dat_dec_inst = d_io_dat_dec_inst; // @[core.scala 28:14]
  assign c_io_dat_exe_br_eq = d_io_dat_exe_br_eq; // @[core.scala 28:14]
  assign c_io_dat_exe_br_lt = d_io_dat_exe_br_lt; // @[core.scala 28:14]
  assign c_io_dat_exe_br_ltu = d_io_dat_exe_br_ltu; // @[core.scala 28:14]
  assign c_io_dat_exe_br_type = d_io_dat_exe_br_type; // @[core.scala 28:14]
  assign c_io_dat_mem_ctrl_dmem_val = d_io_dat_mem_ctrl_dmem_val; // @[core.scala 28:14]
  assign c_io_dat_csr_eret = d_io_dat_csr_eret; // @[core.scala 28:14]
  assign d_clock = clock;
  assign d_reset = reset;
  assign d_io_imem_resp_bits_data = io_imem_resp_bits_data; // @[core.scala 31:12]
  assign d_io_dmem_resp_bits_data = io_dmem_resp_bits_data; // @[core.scala 35:12]
  assign d_io_ctl_dec_stall = c_io_ctl_dec_stall; // @[core.scala 27:14]
  assign d_io_ctl_full_stall = c_io_ctl_full_stall; // @[core.scala 27:14]
  assign d_io_ctl_exe_pc_sel = c_io_ctl_exe_pc_sel; // @[core.scala 27:14]
  assign d_io_ctl_br_type = c_io_ctl_br_type; // @[core.scala 27:14]
  assign d_io_ctl_if_kill = c_io_ctl_if_kill; // @[core.scala 27:14]
  assign d_io_ctl_dec_kill = c_io_ctl_dec_kill; // @[core.scala 27:14]
  assign d_io_ctl_op1_sel = c_io_ctl_op1_sel; // @[core.scala 27:14]
  assign d_io_ctl_op2_sel = c_io_ctl_op2_sel; // @[core.scala 27:14]
  assign d_io_ctl_alu_fun = c_io_ctl_alu_fun; // @[core.scala 27:14]
  assign d_io_ctl_wb_sel = c_io_ctl_wb_sel; // @[core.scala 27:14]
  assign d_io_ctl_rf_wen = c_io_ctl_rf_wen; // @[core.scala 27:14]
  assign d_io_ctl_mem_val = c_io_ctl_mem_val; // @[core.scala 27:14]
  assign d_io_ctl_mem_fcn = c_io_ctl_mem_fcn; // @[core.scala 27:14]
  assign d_io_ctl_mem_typ = c_io_ctl_mem_typ; // @[core.scala 27:14]
  assign d_io_ctl_csr_cmd = c_io_ctl_csr_cmd; // @[core.scala 27:14]
  assign d_io_ctl_fencei = c_io_ctl_fencei; // @[core.scala 27:14]
  assign d_io_ctl_pipeline_kill = c_io_ctl_pipeline_kill; // @[core.scala 27:14]
  assign d_io_ctl_mem_exception = c_io_ctl_mem_exception; // @[core.scala 27:14]
endmodule
module AsyncReadMem(
  input         metaReset,
  input         clock,
  input  [20:0] io_dataInstr_0_addr,
  output [31:0] io_dataInstr_0_data,
  input  [20:0] io_dw_addr,
  input  [31:0] io_dw_data,
  input         io_dw_en
);
  wire  mem_sparse_metaReset; // @[memory.scala 93:28]
  wire  mem_sparse_clock; // @[memory.scala 93:28]
  wire [20:0] mem_sparse_io_w_1_addr; // @[memory.scala 93:28]
  wire  mem_sparse_io_w_1_en; // @[memory.scala 93:28]
  wire [7:0] mem_sparse_io_w_1_data; // @[memory.scala 93:28]
  wire [20:0] mem_sparse_io_r_0_addr; // @[memory.scala 93:28]
  wire [7:0] mem_sparse_io_r_0_data; // @[memory.scala 93:28]
  wire  mem_sparse_0_metaReset; // @[memory.scala 93:28]
  wire  mem_sparse_0_clock; // @[memory.scala 93:28]
  wire [20:0] mem_sparse_0_io_w_1_addr; // @[memory.scala 93:28]
  wire  mem_sparse_0_io_w_1_en; // @[memory.scala 93:28]
  wire [7:0] mem_sparse_0_io_w_1_data; // @[memory.scala 93:28]
  wire [20:0] mem_sparse_0_io_r_0_addr; // @[memory.scala 93:28]
  wire [7:0] mem_sparse_0_io_r_0_data; // @[memory.scala 93:28]
  wire  mem_sparse_1_metaReset; // @[memory.scala 93:28]
  wire  mem_sparse_1_clock; // @[memory.scala 93:28]
  wire [20:0] mem_sparse_1_io_w_1_addr; // @[memory.scala 93:28]
  wire  mem_sparse_1_io_w_1_en; // @[memory.scala 93:28]
  wire [7:0] mem_sparse_1_io_w_1_data; // @[memory.scala 93:28]
  wire [20:0] mem_sparse_1_io_r_0_addr; // @[memory.scala 93:28]
  wire [7:0] mem_sparse_1_io_r_0_data; // @[memory.scala 93:28]
  wire  mem_sparse_2_metaReset; // @[memory.scala 93:28]
  wire  mem_sparse_2_clock; // @[memory.scala 93:28]
  wire [20:0] mem_sparse_2_io_w_1_addr; // @[memory.scala 93:28]
  wire  mem_sparse_2_io_w_1_en; // @[memory.scala 93:28]
  wire [7:0] mem_sparse_2_io_w_1_data; // @[memory.scala 93:28]
  wire [20:0] mem_sparse_2_io_r_0_addr; // @[memory.scala 93:28]
  wire [7:0] mem_sparse_2_io_r_0_data; // @[memory.scala 93:28]
  wire [7:0] underlying_1__T_54_data = mem_sparse_0_io_r_0_data; // @[memory.scala 93:28]
  wire [7:0] underlying_0__T_54_data = mem_sparse_io_r_0_data; // @[memory.scala 93:28]
  wire [15:0] _T_68 = {underlying_1__T_54_data,underlying_0__T_54_data}; // @[memory.scala 82:55]
  wire [7:0] underlying_3__T_54_data = mem_sparse_2_io_r_0_data; // @[memory.scala 93:28]
  wire [7:0] underlying_2__T_54_data = mem_sparse_1_io_r_0_data; // @[memory.scala 93:28]
  wire [15:0] _T_69 = {underlying_3__T_54_data,underlying_2__T_54_data}; // @[memory.scala 82:55]
  SparseMem_0 mem_sparse ( // @[memory.scala 93:28]
    .metaReset(mem_sparse_metaReset),
    .clock(mem_sparse_clock),
    .io_w_1_addr(mem_sparse_io_w_1_addr),
    .io_w_1_en(mem_sparse_io_w_1_en),
    .io_w_1_data(mem_sparse_io_w_1_data),
    .io_r_0_addr(mem_sparse_io_r_0_addr),
    .io_r_0_data(mem_sparse_io_r_0_data)
  );
  SparseMem_0 mem_sparse_0 ( // @[memory.scala 93:28]
    .metaReset(mem_sparse_0_metaReset),
    .clock(mem_sparse_0_clock),
    .io_w_1_addr(mem_sparse_0_io_w_1_addr),
    .io_w_1_en(mem_sparse_0_io_w_1_en),
    .io_w_1_data(mem_sparse_0_io_w_1_data),
    .io_r_0_addr(mem_sparse_0_io_r_0_addr),
    .io_r_0_data(mem_sparse_0_io_r_0_data)
  );
  SparseMem_0 mem_sparse_1 ( // @[memory.scala 93:28]
    .metaReset(mem_sparse_1_metaReset),
    .clock(mem_sparse_1_clock),
    .io_w_1_addr(mem_sparse_1_io_w_1_addr),
    .io_w_1_en(mem_sparse_1_io_w_1_en),
    .io_w_1_data(mem_sparse_1_io_w_1_data),
    .io_r_0_addr(mem_sparse_1_io_r_0_addr),
    .io_r_0_data(mem_sparse_1_io_r_0_data)
  );
  SparseMem_0 mem_sparse_2 ( // @[memory.scala 93:28]
    .metaReset(mem_sparse_2_metaReset),
    .clock(mem_sparse_2_clock),
    .io_w_1_addr(mem_sparse_2_io_w_1_addr),
    .io_w_1_en(mem_sparse_2_io_w_1_en),
    .io_w_1_data(mem_sparse_2_io_w_1_data),
    .io_r_0_addr(mem_sparse_2_io_r_0_addr),
    .io_r_0_data(mem_sparse_2_io_r_0_data)
  );
  assign mem_sparse_metaReset = metaReset;
  assign mem_sparse_0_metaReset = metaReset;
  assign mem_sparse_1_metaReset = metaReset;
  assign mem_sparse_2_metaReset = metaReset;
  assign io_dataInstr_0_data = {_T_69,_T_68}; // @[memory.scala 82:16]
  assign mem_sparse_clock = clock;
  assign mem_sparse_io_w_1_addr = io_dw_addr;
  assign mem_sparse_io_w_1_en = io_dw_en;
  assign mem_sparse_io_w_1_data = io_dw_data[7:0];
  assign mem_sparse_io_r_0_addr = io_dataInstr_0_addr;
  assign mem_sparse_0_clock = clock;
  assign mem_sparse_0_io_w_1_addr = io_dw_addr;
  assign mem_sparse_0_io_w_1_en = io_dw_en;
  assign mem_sparse_0_io_w_1_data = io_dw_data[15:8];
  assign mem_sparse_0_io_r_0_addr = io_dataInstr_0_addr;
  assign mem_sparse_1_clock = clock;
  assign mem_sparse_1_io_w_1_addr = io_dw_addr;
  assign mem_sparse_1_io_w_1_en = io_dw_en;
  assign mem_sparse_1_io_w_1_data = io_dw_data[23:16];
  assign mem_sparse_1_io_r_0_addr = io_dataInstr_0_addr;
  assign mem_sparse_2_clock = clock;
  assign mem_sparse_2_io_w_1_addr = io_dw_addr;
  assign mem_sparse_2_io_w_1_en = io_dw_en;
  assign mem_sparse_2_io_w_1_data = io_dw_data[31:24];
  assign mem_sparse_2_io_r_0_addr = io_dataInstr_0_addr;
endmodule
module SparseMem_0(
  input         metaReset,
  input         clock,
  input  [20:0] io_w_1_addr,
  input         io_w_1_en,
  input  [7:0]  io_w_1_data,
  input  [20:0] io_r_0_addr,
  output [7:0]  io_r_0_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] mem [0:31];
  wire [7:0] mem__T_152_data;
  wire [4:0] mem__T_152_addr;
  wire [7:0] mem__T_274_data;
  wire [4:0] mem__T_274_addr;
  wire [7:0] mem__T_396_data;
  wire [4:0] mem__T_396_addr;
  wire [7:0] mem__T_528_data;
  wire [4:0] mem__T_528_addr;
  wire  mem__T_528_mask;
  wire  mem__T_528_en;
  wire [7:0] mem__T_656_data;
  wire [4:0] mem__T_656_addr;
  wire  mem__T_656_mask;
  wire  mem__T_656_en;
  reg [20:0] addresses_0_bits;
  reg [20:0] addresses_1_bits;
  reg [20:0] addresses_2_bits;
  reg [20:0] addresses_3_bits;
  reg [20:0] addresses_4_bits;
  reg [20:0] addresses_5_bits;
  reg [20:0] addresses_6_bits;
  reg [20:0] addresses_7_bits;
  reg [20:0] addresses_8_bits;
  reg [20:0] addresses_9_bits;
  reg [20:0] addresses_10_bits;
  reg [20:0] addresses_11_bits;
  reg [20:0] addresses_12_bits;
  reg [20:0] addresses_13_bits;
  reg [20:0] addresses_14_bits;
  reg [20:0] addresses_15_bits;
  reg [20:0] addresses_16_bits;
  reg [20:0] addresses_17_bits;
  reg [20:0] addresses_18_bits;
  reg [20:0] addresses_19_bits;
  reg [20:0] addresses_20_bits;
  reg [20:0] addresses_21_bits;
  reg [20:0] addresses_22_bits;
  reg [20:0] addresses_23_bits;
  reg [20:0] addresses_24_bits;
  reg [20:0] addresses_25_bits;
  reg [20:0] addresses_26_bits;
  reg [20:0] addresses_27_bits;
  reg [20:0] addresses_28_bits;
  reg [20:0] addresses_29_bits;
  reg [20:0] addresses_30_bits;
  reg [20:0] addresses_31_bits;
  wire  _T_33 = addresses_0_bits == io_r_0_addr;
  wire  _T_35 = addresses_1_bits == io_r_0_addr;
  wire  _T_37 = addresses_2_bits == io_r_0_addr;
  wire  _T_39 = addresses_3_bits == io_r_0_addr;
  wire  _T_41 = addresses_4_bits == io_r_0_addr;
  wire  _T_43 = addresses_5_bits == io_r_0_addr;
  wire  _T_45 = addresses_6_bits == io_r_0_addr;
  wire  _T_47 = addresses_7_bits == io_r_0_addr;
  wire  _T_49 = addresses_8_bits == io_r_0_addr;
  wire  _T_51 = addresses_9_bits == io_r_0_addr;
  wire  _T_53 = addresses_10_bits == io_r_0_addr;
  wire  _T_55 = addresses_11_bits == io_r_0_addr;
  wire  _T_57 = addresses_12_bits == io_r_0_addr;
  wire  _T_59 = addresses_13_bits == io_r_0_addr;
  wire  _T_61 = addresses_14_bits == io_r_0_addr;
  wire  _T_63 = addresses_15_bits == io_r_0_addr;
  wire  _T_65 = addresses_16_bits == io_r_0_addr;
  wire  _T_67 = addresses_17_bits == io_r_0_addr;
  wire  _T_69 = addresses_18_bits == io_r_0_addr;
  wire  _T_71 = addresses_19_bits == io_r_0_addr;
  wire  _T_73 = addresses_20_bits == io_r_0_addr;
  wire  _T_75 = addresses_21_bits == io_r_0_addr;
  wire  _T_77 = addresses_22_bits == io_r_0_addr;
  wire  _T_79 = addresses_23_bits == io_r_0_addr;
  wire  _T_81 = addresses_24_bits == io_r_0_addr;
  wire  _T_83 = addresses_25_bits == io_r_0_addr;
  wire  _T_85 = addresses_26_bits == io_r_0_addr;
  wire  _T_87 = addresses_27_bits == io_r_0_addr;
  wire  _T_89 = addresses_28_bits == io_r_0_addr;
  wire  _T_91 = addresses_29_bits == io_r_0_addr;
  wire  _T_93 = addresses_30_bits == io_r_0_addr;
  wire  _T_95 = addresses_31_bits == io_r_0_addr;
  wire [7:0] _T_104 = {_T_47,_T_45,_T_43,_T_41,_T_39,_T_37,_T_35,_T_33};
  wire [15:0] _T_112 = {_T_63,_T_61,_T_59,_T_57,_T_55,_T_53,_T_51,_T_49,_T_104};
  wire [7:0] _T_119 = {_T_79,_T_77,_T_75,_T_73,_T_71,_T_69,_T_67,_T_65};
  wire [31:0] _T_128 = {_T_95,_T_93,_T_91,_T_89,_T_87,_T_85,_T_83,_T_81,_T_119,_T_112};
  wire  _T_129 = _T_128 != 32'h0;
  wire  _T_132 = |_T_128[31:16];
  wire [15:0] _T_133 = _T_128[31:16] | _T_128[15:0];
  wire  _T_136 = |_T_133[15:8];
  wire [7:0] _T_137 = _T_133[15:8] | _T_133[7:0];
  wire  _T_140 = |_T_137[7:4];
  wire [3:0] _T_141 = _T_137[7:4] | _T_137[3:0];
  wire  _T_144 = |_T_141[3:2];
  wire [1:0] _T_145 = _T_141[3:2] | _T_141[1:0];
  wire [3:0] _T_149 = {_T_136,_T_140,_T_144,_T_145[1]};
  wire  _T_155 = addresses_0_bits == 21'h0;
  wire  _T_157 = addresses_1_bits == 21'h0;
  wire  _T_159 = addresses_2_bits == 21'h0;
  wire  _T_161 = addresses_3_bits == 21'h0;
  wire  _T_163 = addresses_4_bits == 21'h0;
  wire  _T_165 = addresses_5_bits == 21'h0;
  wire  _T_167 = addresses_6_bits == 21'h0;
  wire  _T_169 = addresses_7_bits == 21'h0;
  wire  _T_171 = addresses_8_bits == 21'h0;
  wire  _T_173 = addresses_9_bits == 21'h0;
  wire  _T_175 = addresses_10_bits == 21'h0;
  wire  _T_177 = addresses_11_bits == 21'h0;
  wire  _T_179 = addresses_12_bits == 21'h0;
  wire  _T_181 = addresses_13_bits == 21'h0;
  wire  _T_183 = addresses_14_bits == 21'h0;
  wire  _T_185 = addresses_15_bits == 21'h0;
  wire  _T_187 = addresses_16_bits == 21'h0;
  wire  _T_189 = addresses_17_bits == 21'h0;
  wire  _T_191 = addresses_18_bits == 21'h0;
  wire  _T_193 = addresses_19_bits == 21'h0;
  wire  _T_195 = addresses_20_bits == 21'h0;
  wire  _T_197 = addresses_21_bits == 21'h0;
  wire  _T_199 = addresses_22_bits == 21'h0;
  wire  _T_201 = addresses_23_bits == 21'h0;
  wire  _T_203 = addresses_24_bits == 21'h0;
  wire  _T_205 = addresses_25_bits == 21'h0;
  wire  _T_207 = addresses_26_bits == 21'h0;
  wire  _T_209 = addresses_27_bits == 21'h0;
  wire  _T_211 = addresses_28_bits == 21'h0;
  wire  _T_213 = addresses_29_bits == 21'h0;
  wire  _T_215 = addresses_30_bits == 21'h0;
  wire  _T_217 = addresses_31_bits == 21'h0;
  wire [7:0] _T_226 = {_T_169,_T_167,_T_165,_T_163,_T_161,_T_159,_T_157,_T_155};
  wire [15:0] _T_234 = {_T_185,_T_183,_T_181,_T_179,_T_177,_T_175,_T_173,_T_171,_T_226};
  wire [7:0] _T_241 = {_T_201,_T_199,_T_197,_T_195,_T_193,_T_191,_T_189,_T_187};
  wire [31:0] _T_250 = {_T_217,_T_215,_T_213,_T_211,_T_209,_T_207,_T_205,_T_203,_T_241,_T_234};
  wire  _T_251 = _T_250 != 32'h0;
  wire  _T_254 = |_T_250[31:16];
  wire [15:0] _T_255 = _T_250[31:16] | _T_250[15:0];
  wire  _T_258 = |_T_255[15:8];
  wire [7:0] _T_259 = _T_255[15:8] | _T_255[7:0];
  wire  _T_262 = |_T_259[7:4];
  wire [3:0] _T_263 = _T_259[7:4] | _T_259[3:0];
  wire  _T_266 = |_T_263[3:2];
  wire [1:0] _T_267 = _T_263[3:2] | _T_263[1:0];
  wire [3:0] _T_271 = {_T_258,_T_262,_T_266,_T_267[1]};
  wire [4:0] _T_272 = {_T_254,_T_258,_T_262,_T_266,_T_267[1]};
  reg [5:0] nextAddr;
  wire [5:0] _T_400 = nextAddr + 6'h1;
  wire [5:0] _T_524 = _T_251 ? {{1'd0}, _T_272} : nextAddr;
  wire  _T_532 = addresses_0_bits == io_w_1_addr;
  wire  _T_534 = addresses_1_bits == io_w_1_addr;
  wire  _T_536 = addresses_2_bits == io_w_1_addr;
  wire  _T_538 = addresses_3_bits == io_w_1_addr;
  wire  _T_540 = addresses_4_bits == io_w_1_addr;
  wire  _T_542 = addresses_5_bits == io_w_1_addr;
  wire  _T_544 = addresses_6_bits == io_w_1_addr;
  wire  _T_546 = addresses_7_bits == io_w_1_addr;
  wire  _T_548 = addresses_8_bits == io_w_1_addr;
  wire  _T_550 = addresses_9_bits == io_w_1_addr;
  wire  _T_552 = addresses_10_bits == io_w_1_addr;
  wire  _T_554 = addresses_11_bits == io_w_1_addr;
  wire  _T_556 = addresses_12_bits == io_w_1_addr;
  wire  _T_558 = addresses_13_bits == io_w_1_addr;
  wire  _T_560 = addresses_14_bits == io_w_1_addr;
  wire  _T_562 = addresses_15_bits == io_w_1_addr;
  wire  _T_564 = addresses_16_bits == io_w_1_addr;
  wire  _T_566 = addresses_17_bits == io_w_1_addr;
  wire  _T_568 = addresses_18_bits == io_w_1_addr;
  wire  _T_570 = addresses_19_bits == io_w_1_addr;
  wire  _T_572 = addresses_20_bits == io_w_1_addr;
  wire  _T_574 = addresses_21_bits == io_w_1_addr;
  wire  _T_576 = addresses_22_bits == io_w_1_addr;
  wire  _T_578 = addresses_23_bits == io_w_1_addr;
  wire  _T_580 = addresses_24_bits == io_w_1_addr;
  wire  _T_582 = addresses_25_bits == io_w_1_addr;
  wire  _T_584 = addresses_26_bits == io_w_1_addr;
  wire  _T_586 = addresses_27_bits == io_w_1_addr;
  wire  _T_588 = addresses_28_bits == io_w_1_addr;
  wire  _T_590 = addresses_29_bits == io_w_1_addr;
  wire  _T_592 = addresses_30_bits == io_w_1_addr;
  wire  _T_594 = addresses_31_bits == io_w_1_addr;
  wire [7:0] _T_603 = {_T_546,_T_544,_T_542,_T_540,_T_538,_T_536,_T_534,_T_532};
  wire [15:0] _T_611 = {_T_562,_T_560,_T_558,_T_556,_T_554,_T_552,_T_550,_T_548,_T_603};
  wire [7:0] _T_618 = {_T_578,_T_576,_T_574,_T_572,_T_570,_T_568,_T_566,_T_564};
  wire [31:0] _T_627 = {_T_594,_T_592,_T_590,_T_588,_T_586,_T_584,_T_582,_T_580,_T_618,_T_611};
  wire  _T_628 = _T_627 != 32'h0;
  wire  _T_631 = |_T_627[31:16];
  wire [15:0] _T_632 = _T_627[31:16] | _T_627[15:0];
  wire  _T_635 = |_T_632[15:8];
  wire [7:0] _T_636 = _T_632[15:8] | _T_632[7:0];
  wire  _T_639 = |_T_636[7:4];
  wire [3:0] _T_640 = _T_636[7:4] | _T_636[3:0];
  wire  _T_643 = |_T_640[3:2];
  wire [1:0] _T_644 = _T_640[3:2] | _T_640[1:0];
  wire [4:0] _T_649 = {_T_631,_T_635,_T_639,_T_643,_T_644[1]};
  wire  _T_650 = ~_T_628;
  wire  _T_651 = io_w_1_en & _T_650;
  wire [5:0] _T_652 = _T_628 ? {{1'd0}, _T_649} : nextAddr;
  wire [5:0] nextAddrUpdate = _T_651 ? _T_400 : nextAddr;
  wire  _T_659 = nextAddrUpdate <= 6'h20;
  wire  _T_662 = ~_T_659;
  assign mem__T_152_addr = {_T_132,_T_149};
  assign mem__T_152_data = mem[mem__T_152_addr];
  assign mem__T_274_addr = {_T_254,_T_271};
  assign mem__T_274_data = mem[mem__T_274_addr];
  assign mem__T_396_addr = {_T_254,_T_271};
  assign mem__T_396_data = mem[mem__T_396_addr];
  assign mem__T_528_data = 8'h0;
  assign mem__T_528_addr = _T_524[4:0];
  assign mem__T_528_mask = 1'h1;
  assign mem__T_528_en = 1'h0;
  assign mem__T_656_data = io_w_1_data;
  assign mem__T_656_addr = _T_652[4:0];
  assign mem__T_656_mask = 1'h1;
  assign mem__T_656_en = io_w_1_en;
  assign io_r_0_data = _T_129 ? mem__T_152_data : 8'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    mem[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  addresses_0_bits = _RAND_1[20:0];
  _RAND_2 = {1{`RANDOM}};
  addresses_1_bits = _RAND_2[20:0];
  _RAND_3 = {1{`RANDOM}};
  addresses_2_bits = _RAND_3[20:0];
  _RAND_4 = {1{`RANDOM}};
  addresses_3_bits = _RAND_4[20:0];
  _RAND_5 = {1{`RANDOM}};
  addresses_4_bits = _RAND_5[20:0];
  _RAND_6 = {1{`RANDOM}};
  addresses_5_bits = _RAND_6[20:0];
  _RAND_7 = {1{`RANDOM}};
  addresses_6_bits = _RAND_7[20:0];
  _RAND_8 = {1{`RANDOM}};
  addresses_7_bits = _RAND_8[20:0];
  _RAND_9 = {1{`RANDOM}};
  addresses_8_bits = _RAND_9[20:0];
  _RAND_10 = {1{`RANDOM}};
  addresses_9_bits = _RAND_10[20:0];
  _RAND_11 = {1{`RANDOM}};
  addresses_10_bits = _RAND_11[20:0];
  _RAND_12 = {1{`RANDOM}};
  addresses_11_bits = _RAND_12[20:0];
  _RAND_13 = {1{`RANDOM}};
  addresses_12_bits = _RAND_13[20:0];
  _RAND_14 = {1{`RANDOM}};
  addresses_13_bits = _RAND_14[20:0];
  _RAND_15 = {1{`RANDOM}};
  addresses_14_bits = _RAND_15[20:0];
  _RAND_16 = {1{`RANDOM}};
  addresses_15_bits = _RAND_16[20:0];
  _RAND_17 = {1{`RANDOM}};
  addresses_16_bits = _RAND_17[20:0];
  _RAND_18 = {1{`RANDOM}};
  addresses_17_bits = _RAND_18[20:0];
  _RAND_19 = {1{`RANDOM}};
  addresses_18_bits = _RAND_19[20:0];
  _RAND_20 = {1{`RANDOM}};
  addresses_19_bits = _RAND_20[20:0];
  _RAND_21 = {1{`RANDOM}};
  addresses_20_bits = _RAND_21[20:0];
  _RAND_22 = {1{`RANDOM}};
  addresses_21_bits = _RAND_22[20:0];
  _RAND_23 = {1{`RANDOM}};
  addresses_22_bits = _RAND_23[20:0];
  _RAND_24 = {1{`RANDOM}};
  addresses_23_bits = _RAND_24[20:0];
  _RAND_25 = {1{`RANDOM}};
  addresses_24_bits = _RAND_25[20:0];
  _RAND_26 = {1{`RANDOM}};
  addresses_25_bits = _RAND_26[20:0];
  _RAND_27 = {1{`RANDOM}};
  addresses_26_bits = _RAND_27[20:0];
  _RAND_28 = {1{`RANDOM}};
  addresses_27_bits = _RAND_28[20:0];
  _RAND_29 = {1{`RANDOM}};
  addresses_28_bits = _RAND_29[20:0];
  _RAND_30 = {1{`RANDOM}};
  addresses_29_bits = _RAND_30[20:0];
  _RAND_31 = {1{`RANDOM}};
  addresses_30_bits = _RAND_31[20:0];
  _RAND_32 = {1{`RANDOM}};
  addresses_31_bits = _RAND_32[20:0];
  _RAND_33 = {1{`RANDOM}};
  nextAddr = _RAND_33[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_528_en & mem__T_528_mask) begin
      mem[mem__T_528_addr] <= mem__T_528_data;
    end
    if(mem__T_656_en & mem__T_656_mask) begin
      mem[mem__T_656_addr] <= mem__T_656_data;
    end
    if (metaReset) begin
      addresses_0_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h0 == _T_652[4:0]) begin
        addresses_0_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_1_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h1 == _T_652[4:0]) begin
        addresses_1_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_2_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h2 == _T_652[4:0]) begin
        addresses_2_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_3_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h3 == _T_652[4:0]) begin
        addresses_3_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_4_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h4 == _T_652[4:0]) begin
        addresses_4_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_5_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h5 == _T_652[4:0]) begin
        addresses_5_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_6_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h6 == _T_652[4:0]) begin
        addresses_6_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_7_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h7 == _T_652[4:0]) begin
        addresses_7_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_8_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h8 == _T_652[4:0]) begin
        addresses_8_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_9_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h9 == _T_652[4:0]) begin
        addresses_9_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_10_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'ha == _T_652[4:0]) begin
        addresses_10_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_11_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'hb == _T_652[4:0]) begin
        addresses_11_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_12_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'hc == _T_652[4:0]) begin
        addresses_12_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_13_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'hd == _T_652[4:0]) begin
        addresses_13_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_14_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'he == _T_652[4:0]) begin
        addresses_14_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_15_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'hf == _T_652[4:0]) begin
        addresses_15_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_16_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h10 == _T_652[4:0]) begin
        addresses_16_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_17_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h11 == _T_652[4:0]) begin
        addresses_17_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_18_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h12 == _T_652[4:0]) begin
        addresses_18_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_19_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h13 == _T_652[4:0]) begin
        addresses_19_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_20_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h14 == _T_652[4:0]) begin
        addresses_20_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_21_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h15 == _T_652[4:0]) begin
        addresses_21_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_22_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h16 == _T_652[4:0]) begin
        addresses_22_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_23_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h17 == _T_652[4:0]) begin
        addresses_23_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_24_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h18 == _T_652[4:0]) begin
        addresses_24_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_25_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h19 == _T_652[4:0]) begin
        addresses_25_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_26_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h1a == _T_652[4:0]) begin
        addresses_26_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_27_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h1b == _T_652[4:0]) begin
        addresses_27_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_28_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h1c == _T_652[4:0]) begin
        addresses_28_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_29_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h1d == _T_652[4:0]) begin
        addresses_29_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_30_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h1e == _T_652[4:0]) begin
        addresses_30_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_31_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h1f == _T_652[4:0]) begin
        addresses_31_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      nextAddr <= 6'h0;
    end else if (_T_651) begin
      nextAddr <= _T_400;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif

    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif

    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AsyncScratchPadMemory(
  input         metaReset,
  input         clock,
  input         io_core_ports_0_req_valid,
  input  [31:0] io_core_ports_0_req_bits_addr,
  input  [31:0] io_core_ports_0_req_bits_data,
  input         io_core_ports_0_req_bits_fcn,
  input  [2:0]  io_core_ports_0_req_bits_typ,
  output        io_core_ports_0_resp_valid,
  output [31:0] io_core_ports_0_resp_bits_data,
  output        _GEN_4_0,
  output        _GEN_1_1,
  output        _GEN_0_1,
  output        _GEN_3_1,
  output        _GEN_5_0,
  output        _GEN_2_0
);
  wire  async_data_metaReset; // @[memory.scala 137:27]
  wire  async_data_clock; // @[memory.scala 137:27]
  wire [20:0] async_data_io_dataInstr_0_addr; // @[memory.scala 137:27]
  wire [31:0] async_data_io_dataInstr_0_data; // @[memory.scala 137:27]
  wire [20:0] async_data_io_dw_addr; // @[memory.scala 137:27]
  wire [31:0] async_data_io_dw_data; // @[memory.scala 137:27]
  wire  async_data_io_dw_en; // @[memory.scala 137:27]
  wire  _T_230 = io_core_ports_0_req_bits_typ == 3'h1; // @[memory.scala 153:17]
  wire [23:0] _T_235 = async_data_io_dataInstr_0_data[7] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_237 = {_T_235,async_data_io_dataInstr_0_data[7:0]}; // @[Cat.scala 30:58]
  wire  _T_238 = io_core_ports_0_req_bits_typ == 3'h2; // @[memory.scala 154:17]
  wire [15:0] _T_243 = async_data_io_dataInstr_0_data[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_245 = {_T_243,async_data_io_dataInstr_0_data[15:0]}; // @[Cat.scala 30:58]
  wire  _T_246 = io_core_ports_0_req_bits_typ == 3'h5; // @[memory.scala 155:17]
  wire [31:0] _T_253 = {24'h0,async_data_io_dataInstr_0_data[7:0]}; // @[Cat.scala 30:58]
  wire  _T_254 = io_core_ports_0_req_bits_typ == 3'h6; // @[memory.scala 156:17]
  wire [31:0] _T_261 = {16'h0,async_data_io_dataInstr_0_data[15:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_262 = _T_254 ? _T_261 : async_data_io_dataInstr_0_data; // @[Mux.scala 61:16]
  wire [31:0] _T_263 = _T_246 ? _T_253 : _T_262; // @[Mux.scala 61:16]
  wire [31:0] _T_264 = _T_238 ? _T_245 : _T_263; // @[Mux.scala 61:16]
  wire [4:0] _T_273 = {io_core_ports_0_req_bits_addr[1:0], 3'h0}; // @[memory.scala 161:86]
  wire [62:0] _GEN_8 = {{31'd0}, io_core_ports_0_req_bits_data}; // @[memory.scala 161:67]
  wire [62:0] _T_274 = _GEN_8 << _T_273; // @[memory.scala 161:67]
  wire [31:0] _T_277 = {io_core_ports_0_req_bits_addr[31:2],2'h0}; // @[Cat.scala 30:58]
  AsyncReadMem async_data ( // @[memory.scala 137:27]
    .metaReset(async_data_metaReset),
    .clock(async_data_clock),
    .io_dataInstr_0_addr(async_data_io_dataInstr_0_addr),
    .io_dataInstr_0_data(async_data_io_dataInstr_0_data),
    .io_dw_addr(async_data_io_dw_addr),
    .io_dw_data(async_data_io_dw_data),
    .io_dw_en(async_data_io_dw_en)
  );
  assign async_data_metaReset = metaReset;
  assign io_core_ports_0_resp_valid = io_core_ports_0_req_valid; // @[memory.scala 142:35]
  assign io_core_ports_0_resp_bits_data = _T_230 ? _T_237 : _T_264; // @[memory.scala 152:40]
  assign _GEN_4_0 = io_core_ports_0_req_bits_typ == 3'h2;
  assign _GEN_1_1 = async_data_io_dataInstr_0_data[15];
  assign _GEN_0_1 = async_data_io_dataInstr_0_data[7];
  assign _GEN_3_1 = io_core_ports_0_req_bits_typ == 3'h5;
  assign _GEN_5_0 = io_core_ports_0_req_bits_typ == 3'h1;
  assign _GEN_2_0 = io_core_ports_0_req_bits_typ == 3'h6;
  assign async_data_clock = clock;
  assign async_data_io_dataInstr_0_addr = io_core_ports_0_req_bits_addr[20:0]; // @[memory.scala 144:39]
  assign async_data_io_dw_addr = _T_277[20:0]; // @[memory.scala 162:29]
  assign async_data_io_dw_data = _T_274[31:0]; // @[memory.scala 161:29]
  assign async_data_io_dw_en = io_core_ports_0_req_bits_fcn; // @[memory.scala 158:24]
endmodule
