module ibex_decoder( // @[ibex_decoder.v:1.1-458.10:ibex_decoder.fir@2.2]
  output        branch_in_dec_o, // @[ibex_decoder.v:82.13-82.28:ibex_decoder.fir@3.4]
  output        jump_in_dec_o, // @[ibex_decoder.v:81.13-81.26:ibex_decoder.fir@4.4]
  output        data_sign_extension_o, // @[ibex_decoder.v:80.13-80.34:ibex_decoder.fir@5.4]
  output [1:0]  data_type_o, // @[ibex_decoder.v:79.19-79.30:ibex_decoder.fir@6.4]
  output        data_we_o, // @[ibex_decoder.v:78.13-78.22:ibex_decoder.fir@7.4]
  output        data_req_o, // @[ibex_decoder.v:77.13-77.23:ibex_decoder.fir@8.4]
  output        csr_pipe_flush_o, // @[ibex_decoder.v:76.13-76.29:ibex_decoder.fir@9.4]
  output [1:0]  csr_op_o, // @[ibex_decoder.v:75.19-75.27:ibex_decoder.fir@10.4]
  output        csr_access_o, // @[ibex_decoder.v:74.13-74.25:ibex_decoder.fir@11.4]
  output [1:0]  multdiv_signed_mode_o, // @[ibex_decoder.v:73.19-73.40:ibex_decoder.fir@12.4]
  output [1:0]  multdiv_operator_o, // @[ibex_decoder.v:72.19-72.37:ibex_decoder.fir@13.4]
  output        div_en_o, // @[ibex_decoder.v:71.13-71.21:ibex_decoder.fir@14.4]
  output        mult_en_o, // @[ibex_decoder.v:70.13-70.22:ibex_decoder.fir@15.4]
  output        alu_op_b_mux_sel_o, // @[ibex_decoder.v:69.13-69.31:ibex_decoder.fir@16.4]
  output [1:0]  alu_op_a_mux_sel_o, // @[ibex_decoder.v:68.19-68.37:ibex_decoder.fir@17.4]
  output [4:0]  alu_operator_o, // @[ibex_decoder.v:67.19-67.33:ibex_decoder.fir@18.4]
  output [4:0]  regfile_waddr_o, // @[ibex_decoder.v:66.20-66.35:ibex_decoder.fir@19.4]
  output [4:0]  regfile_raddr_b_o, // @[ibex_decoder.v:65.20-65.37:ibex_decoder.fir@20.4]
  output [4:0]  regfile_raddr_a_o, // @[ibex_decoder.v:64.20-64.37:ibex_decoder.fir@21.4]
  output        regfile_we_o, // @[ibex_decoder.v:63.14-63.26:ibex_decoder.fir@22.4]
  output [1:0]  regfile_wdata_sel_o, // @[ibex_decoder.v:62.19-62.38:ibex_decoder.fir@23.4]
  output [31:0] zimm_rs1_type_o, // @[ibex_decoder.v:61.21-61.36:ibex_decoder.fir@24.4]
  output [31:0] imm_j_type_o, // @[ibex_decoder.v:60.21-60.33:ibex_decoder.fir@25.4]
  output [31:0] imm_u_type_o, // @[ibex_decoder.v:59.21-59.33:ibex_decoder.fir@26.4]
  output [31:0] imm_b_type_o, // @[ibex_decoder.v:58.21-58.33:ibex_decoder.fir@27.4]
  output [31:0] imm_s_type_o, // @[ibex_decoder.v:57.21-57.33:ibex_decoder.fir@28.4]
  output [31:0] imm_i_type_o, // @[ibex_decoder.v:56.21-56.33:ibex_decoder.fir@29.4]
  output [2:0]  imm_b_mux_sel_o, // @[ibex_decoder.v:55.19-55.34:ibex_decoder.fir@30.4]
  output        imm_a_mux_sel_o, // @[ibex_decoder.v:54.13-54.28:ibex_decoder.fir@31.4]
  input         illegal_c_insn_i, // @[ibex_decoder.v:53.13-53.29:ibex_decoder.fir@32.4]
  input  [31:0] instr_rdata_i, // @[ibex_decoder.v:52.20-52.33:ibex_decoder.fir@33.4]
  input         instr_new_i, // @[ibex_decoder.v:51.13-51.24:ibex_decoder.fir@34.4]
  output        jump_set_o, // @[ibex_decoder.v:50.13-50.23:ibex_decoder.fir@35.4]
  output        wfi_insn_o, // @[ibex_decoder.v:49.13-49.23:ibex_decoder.fir@36.4]
  output        ecall_insn_o, // @[ibex_decoder.v:48.13-48.25:ibex_decoder.fir@37.4]
  output        dret_insn_o, // @[ibex_decoder.v:47.13-47.24:ibex_decoder.fir@38.4]
  output        mret_insn_o, // @[ibex_decoder.v:46.13-46.24:ibex_decoder.fir@39.4]
  output        ebrk_insn_o, // @[ibex_decoder.v:45.13-45.24:ibex_decoder.fir@40.4]
  output        illegal_insn_o // @[ibex_decoder.v:44.14-44.28:ibex_decoder.fir@41.4]
);
  wire [4:0] _GEN_0; // @[ibex_decoder.v:406.12-406.32:ibex_decoder.fir@292.4]
  wire [4:0] _GEN_1; // @[ibex_decoder.v:406.38-406.58:ibex_decoder.fir@291.4]
  wire [6:0] _GEN_4; // @[ibex_decoder.v:290.17-290.44:ibex_decoder.fir@294.4]
  wire [11:0] _GEN_10; // @[ibex_decoder.v:121.12-121.53:ibex_decoder.fir@306.4]
  wire  _GEN_24; // @[:ibex_decoder.fir@324.4]
  wire [12:0] _GEN_27; // @[:ibex_decoder.fir@324.4]
  wire [13:0] _GEN_29; // @[:ibex_decoder.fir@324.4]
  wire [14:0] _GEN_31; // @[:ibex_decoder.fir@324.4]
  wire [15:0] _GEN_33; // @[:ibex_decoder.fir@324.4]
  wire [16:0] _GEN_35; // @[:ibex_decoder.fir@324.4]
  wire [17:0] _GEN_37; // @[:ibex_decoder.fir@324.4]
  wire [18:0] _GEN_39; // @[:ibex_decoder.fir@324.4]
  wire [19:0] _GEN_41; // @[:ibex_decoder.fir@324.4]
  wire [20:0] _GEN_43; // @[:ibex_decoder.fir@324.4]
  wire [21:0] _GEN_45; // @[:ibex_decoder.fir@324.4]
  wire [22:0] _GEN_47; // @[:ibex_decoder.fir@324.4]
  wire [23:0] _GEN_49; // @[:ibex_decoder.fir@324.4]
  wire [24:0] _GEN_51; // @[:ibex_decoder.fir@324.4]
  wire [25:0] _GEN_53; // @[:ibex_decoder.fir@324.4]
  wire [26:0] _GEN_55; // @[:ibex_decoder.fir@324.4]
  wire [27:0] _GEN_57; // @[:ibex_decoder.fir@324.4]
  wire [28:0] _GEN_59; // @[:ibex_decoder.fir@324.4]
  wire [29:0] _GEN_61; // @[:ibex_decoder.fir@324.4]
  wire [30:0] _GEN_63; // @[:ibex_decoder.fir@324.4]
  wire [11:0] _GEN_67; // @[:ibex_decoder.fir@325.4]
  wire [12:0] _GEN_69; // @[:ibex_decoder.fir@325.4]
  wire [13:0] _GEN_71; // @[:ibex_decoder.fir@325.4]
  wire [14:0] _GEN_73; // @[:ibex_decoder.fir@325.4]
  wire [15:0] _GEN_75; // @[:ibex_decoder.fir@325.4]
  wire [16:0] _GEN_77; // @[:ibex_decoder.fir@325.4]
  wire [17:0] _GEN_79; // @[:ibex_decoder.fir@325.4]
  wire [18:0] _GEN_81; // @[:ibex_decoder.fir@325.4]
  wire [19:0] _GEN_83; // @[:ibex_decoder.fir@325.4]
  wire [20:0] _GEN_85; // @[:ibex_decoder.fir@325.4]
  wire [21:0] _GEN_87; // @[:ibex_decoder.fir@325.4]
  wire [22:0] _GEN_89; // @[:ibex_decoder.fir@325.4]
  wire [23:0] _GEN_91; // @[:ibex_decoder.fir@325.4]
  wire [24:0] _GEN_93; // @[:ibex_decoder.fir@325.4]
  wire [25:0] _GEN_95; // @[:ibex_decoder.fir@325.4]
  wire [26:0] _GEN_97; // @[:ibex_decoder.fir@325.4]
  wire [27:0] _GEN_99; // @[:ibex_decoder.fir@325.4]
  wire [28:0] _GEN_101; // @[:ibex_decoder.fir@325.4]
  wire [29:0] _GEN_103; // @[:ibex_decoder.fir@325.4]
  wire [30:0] _GEN_105; // @[:ibex_decoder.fir@325.4]
  wire [3:0] _GEN_106; // @[:ibex_decoder.fir@326.4]
  wire [5:0] _GEN_107; // @[:ibex_decoder.fir@326.4]
  wire [4:0] _GEN_108; // @[:ibex_decoder.fir@326.4]
  wire  _GEN_109; // @[:ibex_decoder.fir@326.4]
  wire [10:0] _GEN_110; // @[:ibex_decoder.fir@326.4]
  wire [11:0] _GEN_112; // @[:ibex_decoder.fir@326.4]
  wire [12:0] _GEN_114; // @[:ibex_decoder.fir@326.4]
  wire [13:0] _GEN_116; // @[:ibex_decoder.fir@326.4]
  wire [14:0] _GEN_118; // @[:ibex_decoder.fir@326.4]
  wire [15:0] _GEN_120; // @[:ibex_decoder.fir@326.4]
  wire [16:0] _GEN_122; // @[:ibex_decoder.fir@326.4]
  wire [17:0] _GEN_124; // @[:ibex_decoder.fir@326.4]
  wire [18:0] _GEN_126; // @[:ibex_decoder.fir@326.4]
  wire [19:0] _GEN_128; // @[:ibex_decoder.fir@326.4]
  wire [20:0] _GEN_130; // @[:ibex_decoder.fir@326.4]
  wire [21:0] _GEN_132; // @[:ibex_decoder.fir@326.4]
  wire [22:0] _GEN_134; // @[:ibex_decoder.fir@326.4]
  wire [23:0] _GEN_136; // @[:ibex_decoder.fir@326.4]
  wire [24:0] _GEN_138; // @[:ibex_decoder.fir@326.4]
  wire [25:0] _GEN_140; // @[:ibex_decoder.fir@326.4]
  wire [26:0] _GEN_142; // @[:ibex_decoder.fir@326.4]
  wire [27:0] _GEN_144; // @[:ibex_decoder.fir@326.4]
  wire [28:0] _GEN_146; // @[:ibex_decoder.fir@326.4]
  wire [29:0] _GEN_148; // @[:ibex_decoder.fir@326.4]
  wire [30:0] _GEN_150; // @[:ibex_decoder.fir@326.4]
  wire [19:0] _GEN_151; // @[:ibex_decoder.fir@327.4]
  wire [9:0] _GEN_152; // @[:ibex_decoder.fir@328.4]
  wire  _GEN_153; // @[:ibex_decoder.fir@328.4]
  wire [10:0] _GEN_154; // @[:ibex_decoder.fir@328.4]
  wire [7:0] _GEN_155; // @[:ibex_decoder.fir@328.4]
  wire [11:0] _GEN_156; // @[:ibex_decoder.fir@328.4]
  wire [19:0] _GEN_158; // @[:ibex_decoder.fir@328.4]
  wire [20:0] _GEN_160; // @[:ibex_decoder.fir@328.4]
  wire [21:0] _GEN_162; // @[:ibex_decoder.fir@328.4]
  wire [22:0] _GEN_164; // @[:ibex_decoder.fir@328.4]
  wire [23:0] _GEN_166; // @[:ibex_decoder.fir@328.4]
  wire [24:0] _GEN_168; // @[:ibex_decoder.fir@328.4]
  wire [25:0] _GEN_170; // @[:ibex_decoder.fir@328.4]
  wire [26:0] _GEN_172; // @[:ibex_decoder.fir@328.4]
  wire [27:0] _GEN_174; // @[:ibex_decoder.fir@328.4]
  wire [28:0] _GEN_176; // @[:ibex_decoder.fir@328.4]
  wire [29:0] _GEN_178; // @[:ibex_decoder.fir@328.4]
  wire [30:0] _GEN_180; // @[:ibex_decoder.fir@328.4]
  assign _GEN_0 = instr_rdata_i[19:15]; // @[ibex_decoder.v:406.12-406.32:ibex_decoder.fir@292.4]
  assign _GEN_1 = instr_rdata_i[11:7]; // @[ibex_decoder.v:406.38-406.58:ibex_decoder.fir@291.4]
  assign _GEN_4 = instr_rdata_i[31:25]; // @[ibex_decoder.v:290.17-290.44:ibex_decoder.fir@294.4]
  assign _GEN_10 = instr_rdata_i[31:20]; // @[ibex_decoder.v:121.12-121.53:ibex_decoder.fir@306.4]
  assign _GEN_24 = instr_rdata_i[31]; // @[:ibex_decoder.fir@324.4]
  assign _GEN_27 = {_GEN_24,_GEN_10}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_29 = {_GEN_24,_GEN_27}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_31 = {_GEN_24,_GEN_29}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_33 = {_GEN_24,_GEN_31}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_35 = {_GEN_24,_GEN_33}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_37 = {_GEN_24,_GEN_35}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_39 = {_GEN_24,_GEN_37}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_41 = {_GEN_24,_GEN_39}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_43 = {_GEN_24,_GEN_41}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_45 = {_GEN_24,_GEN_43}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_47 = {_GEN_24,_GEN_45}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_49 = {_GEN_24,_GEN_47}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_51 = {_GEN_24,_GEN_49}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_53 = {_GEN_24,_GEN_51}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_55 = {_GEN_24,_GEN_53}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_57 = {_GEN_24,_GEN_55}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_59 = {_GEN_24,_GEN_57}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_61 = {_GEN_24,_GEN_59}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_63 = {_GEN_24,_GEN_61}; // @[:ibex_decoder.fir@324.4]
  assign _GEN_67 = {_GEN_4,_GEN_1}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_69 = {_GEN_24,_GEN_67}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_71 = {_GEN_24,_GEN_69}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_73 = {_GEN_24,_GEN_71}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_75 = {_GEN_24,_GEN_73}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_77 = {_GEN_24,_GEN_75}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_79 = {_GEN_24,_GEN_77}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_81 = {_GEN_24,_GEN_79}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_83 = {_GEN_24,_GEN_81}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_85 = {_GEN_24,_GEN_83}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_87 = {_GEN_24,_GEN_85}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_89 = {_GEN_24,_GEN_87}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_91 = {_GEN_24,_GEN_89}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_93 = {_GEN_24,_GEN_91}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_95 = {_GEN_24,_GEN_93}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_97 = {_GEN_24,_GEN_95}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_99 = {_GEN_24,_GEN_97}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_101 = {_GEN_24,_GEN_99}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_103 = {_GEN_24,_GEN_101}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_105 = {_GEN_24,_GEN_103}; // @[:ibex_decoder.fir@325.4]
  assign _GEN_106 = instr_rdata_i[11:8]; // @[:ibex_decoder.fir@326.4]
  assign _GEN_107 = instr_rdata_i[30:25]; // @[:ibex_decoder.fir@326.4]
  assign _GEN_108 = {_GEN_106,1'h0}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_109 = instr_rdata_i[7]; // @[:ibex_decoder.fir@326.4]
  assign _GEN_110 = {_GEN_107,_GEN_108}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_112 = {_GEN_109,_GEN_110}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_114 = {_GEN_24,_GEN_112}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_116 = {_GEN_24,_GEN_114}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_118 = {_GEN_24,_GEN_116}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_120 = {_GEN_24,_GEN_118}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_122 = {_GEN_24,_GEN_120}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_124 = {_GEN_24,_GEN_122}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_126 = {_GEN_24,_GEN_124}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_128 = {_GEN_24,_GEN_126}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_130 = {_GEN_24,_GEN_128}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_132 = {_GEN_24,_GEN_130}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_134 = {_GEN_24,_GEN_132}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_136 = {_GEN_24,_GEN_134}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_138 = {_GEN_24,_GEN_136}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_140 = {_GEN_24,_GEN_138}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_142 = {_GEN_24,_GEN_140}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_144 = {_GEN_24,_GEN_142}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_146 = {_GEN_24,_GEN_144}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_148 = {_GEN_24,_GEN_146}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_150 = {_GEN_24,_GEN_148}; // @[:ibex_decoder.fir@326.4]
  assign _GEN_151 = instr_rdata_i[31:12]; // @[:ibex_decoder.fir@327.4]
  assign _GEN_152 = instr_rdata_i[30:21]; // @[:ibex_decoder.fir@328.4]
  assign _GEN_153 = instr_rdata_i[20]; // @[:ibex_decoder.fir@328.4]
  assign _GEN_154 = {_GEN_152,1'h0}; // @[:ibex_decoder.fir@328.4]
  assign _GEN_155 = instr_rdata_i[19:12]; // @[:ibex_decoder.fir@328.4]
  assign _GEN_156 = {_GEN_153,_GEN_154}; // @[:ibex_decoder.fir@328.4]
  assign _GEN_158 = {_GEN_155,_GEN_156}; // @[:ibex_decoder.fir@328.4]
  assign _GEN_160 = {_GEN_24,_GEN_158}; // @[:ibex_decoder.fir@328.4]
  assign _GEN_162 = {_GEN_24,_GEN_160}; // @[:ibex_decoder.fir@328.4]
  assign _GEN_164 = {_GEN_24,_GEN_162}; // @[:ibex_decoder.fir@328.4]
  assign _GEN_166 = {_GEN_24,_GEN_164}; // @[:ibex_decoder.fir@328.4]
  assign _GEN_168 = {_GEN_24,_GEN_166}; // @[:ibex_decoder.fir@328.4]
  assign _GEN_170 = {_GEN_24,_GEN_168}; // @[:ibex_decoder.fir@328.4]
  assign _GEN_172 = {_GEN_24,_GEN_170}; // @[:ibex_decoder.fir@328.4]
  assign _GEN_174 = {_GEN_24,_GEN_172}; // @[:ibex_decoder.fir@328.4]
  assign _GEN_176 = {_GEN_24,_GEN_174}; // @[:ibex_decoder.fir@328.4]
  assign _GEN_178 = {_GEN_24,_GEN_176}; // @[:ibex_decoder.fir@328.4]
  assign _GEN_180 = {_GEN_24,_GEN_178}; // @[:ibex_decoder.fir@328.4]
  assign branch_in_dec_o = 1'h0;
  assign jump_in_dec_o = 1'h0;
  assign data_sign_extension_o = 1'h0;
  assign data_type_o = 2'h0;
  assign data_we_o = 1'h0;
  assign data_req_o = 1'h0;
  assign csr_pipe_flush_o = 1'h0;
  assign csr_op_o = 2'h0;
  assign csr_access_o = 1'h0;
  assign multdiv_signed_mode_o = 2'h0;
  assign multdiv_operator_o = 2'h0;
  assign div_en_o = 1'h0;
  assign mult_en_o = 1'h0;
  assign alu_op_b_mux_sel_o = 1'h0;
  assign alu_op_a_mux_sel_o = 2'h0;
  assign alu_operator_o = 5'h0;
  assign regfile_waddr_o = instr_rdata_i[11:7];
  assign regfile_raddr_b_o = instr_rdata_i[24:20];
  assign regfile_raddr_a_o = instr_rdata_i[19:15];
  assign regfile_we_o = 1'h0;
  assign regfile_wdata_sel_o = 2'h0;
  assign zimm_rs1_type_o = {27'h0,_GEN_0};
  assign imm_j_type_o = {_GEN_24,_GEN_180};
  assign imm_u_type_o = {_GEN_151,12'h0};
  assign imm_b_type_o = {_GEN_24,_GEN_150};
  assign imm_s_type_o = {_GEN_24,_GEN_105};
  assign imm_i_type_o = {_GEN_24,_GEN_63};
  assign imm_b_mux_sel_o = 3'h0;
  assign imm_a_mux_sel_o = 1'h0;
  assign jump_set_o = 1'h0;
  assign wfi_insn_o = 1'h0;
  assign ecall_insn_o = 1'h0;
  assign dret_insn_o = 1'h0;
  assign mret_insn_o = 1'h0;
  assign ebrk_insn_o = 1'h0;
  assign illegal_insn_o = 1'h0;
endmodule
